
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.bm100_pkg.all;                 -- character ROM type


entity charrom2 is
    port
    (
        clk         : in  std_logic;
        --
        addr_char_i : in  std_logic_vector(7 downto 0);
        addr_line_i : in  std_logic_vector(2 downto 0);
        --
        data_o      : out std_logic_vector(7 downto 0)
    );
end entity charrom2;


architecture rtl of charrom2 is

--  constant rom_init_file : string := "../ROMs/ibm_zg+din.bin";
    constant rom_init_file : string := "../ROMs/zg_m_uml_+inv.bin";

    -- function work with ModelSim (and Xilinx ISE) but not with Quartus 13.1!
    impure function init_crom( filename : string) return T_BM100_MEM is
        type charfile is file of character;
        file data_file  : charfile;
        variable rom    : T_BM100_MEM;
        variable c      : character;
    begin
        if filename'length = 0 then
            report init_crom'instance_name & " no filename given, ROM empty" severity warning;
            return rom;
        end if;

        file_open( data_file, filename, read_mode);
        for index in rom'range loop
            read( data_file, c);
            rom( index) := character'pos( c);
        end loop;
        file_close( data_file);

        return rom;
    end function init_crom;

    --signal crom_array : T_BM100_MEM := init_crom( rom_init_file);

    -- workaround for Quartus
    constant charrom2_init : T_BM100_MEM := (
		16#00#, 16#44#, 16#aa#, 16#aa#, 16#aa#, 16#aa#, 16#44#, 16#00#, -- 0
		16#40#, 16#a0#, 16#0c#, 16#12#, 16#1e#, 16#12#, 16#12#, 16#00#, -- 1
		16#40#, 16#a0#, 16#1c#, 16#12#, 16#1c#, 16#12#, 16#1c#, 16#00#, -- 2
		16#40#, 16#a0#, 16#0c#, 16#12#, 16#10#, 16#12#, 16#0c#, 16#00#, -- 3
		16#40#, 16#a0#, 16#1c#, 16#12#, 16#12#, 16#12#, 16#1c#, 16#00#, -- 4
		16#40#, 16#a0#, 16#1e#, 16#10#, 16#1c#, 16#10#, 16#1e#, 16#00#, -- 5
		16#40#, 16#a0#, 16#1e#, 16#10#, 16#1c#, 16#10#, 16#10#, 16#00#, -- 6
		16#40#, 16#a0#, 16#0c#, 16#12#, 16#10#, 16#16#, 16#0e#, 16#00#, -- 7
		16#40#, 16#a0#, 16#12#, 16#12#, 16#1e#, 16#12#, 16#12#, 16#00#, -- 8
		16#40#, 16#a0#, 16#0e#, 16#04#, 16#04#, 16#04#, 16#0e#, 16#00#, -- 9
		16#00#, 16#00#, 16#8e#, 16#88#, 16#8c#, 16#88#, 16#e8#, 16#00#, -- 10
		16#40#, 16#a0#, 16#12#, 16#14#, 16#18#, 16#14#, 16#12#, 16#00#, -- 11
		16#40#, 16#a0#, 16#10#, 16#10#, 16#10#, 16#10#, 16#1e#, 16#00#, -- 12
		16#00#, 16#00#, 16#6c#, 16#8a#, 16#8c#, 16#8a#, 16#6a#, 16#00#, -- 13
		16#40#, 16#a0#, 16#12#, 16#1a#, 16#16#, 16#12#, 16#12#, 16#00#, -- 14
		16#40#, 16#a0#, 16#0c#, 16#12#, 16#12#, 16#12#, 16#0c#, 16#00#, -- 15
		16#40#, 16#a0#, 16#1c#, 16#12#, 16#1c#, 16#10#, 16#10#, 16#00#, -- 16
		16#40#, 16#a0#, 16#0c#, 16#12#, 16#12#, 16#14#, 16#0a#, 16#00#, -- 17
		16#40#, 16#a0#, 16#1c#, 16#12#, 16#1c#, 16#14#, 16#12#, 16#00#, -- 18
		16#40#, 16#a0#, 16#0e#, 16#10#, 16#0c#, 16#02#, 16#1c#, 16#00#, -- 19
		16#40#, 16#a0#, 16#0e#, 16#04#, 16#04#, 16#04#, 16#04#, 16#00#, -- 20
		16#40#, 16#a0#, 16#12#, 16#12#, 16#12#, 16#12#, 16#0c#, 16#00#, -- 21
		16#40#, 16#a0#, 16#11#, 16#11#, 16#11#, 16#0a#, 16#04#, 16#00#, -- 22
		16#40#, 16#a0#, 16#11#, 16#15#, 16#15#, 16#1b#, 16#11#, 16#00#, -- 23
		16#40#, 16#a0#, 16#11#, 16#0a#, 16#04#, 16#0a#, 16#11#, 16#00#, -- 24
		16#40#, 16#a0#, 16#11#, 16#11#, 16#0a#, 16#04#, 16#04#, 16#00#, -- 25
		16#40#, 16#a0#, 16#1e#, 16#02#, 16#04#, 16#08#, 16#1e#, 16#00#, -- 26
		16#00#, 16#00#, 16#db#, 16#92#, 16#ca#, 16#8a#, 16#db#, 16#00#, -- 27
		16#48#, 16#a8#, 16#08#, 16#08#, 16#08#, 16#08#, 16#08#, 16#00#, -- 28
		16#40#, 16#a0#, 16#0c#, 16#04#, 16#06#, 16#04#, 16#0c#, 16#00#, -- 29
		16#00#, 16#00#, 16#94#, 16#d4#, 16#b4#, 16#94#, 16#96#, 16#00#, -- 30
		16#00#, 16#00#, 16#2e#, 16#68#, 16#2c#, 16#28#, 16#28#, 16#00#, -- 31
		16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, -- 32
		16#10#, 16#10#, 16#10#, 16#10#, 16#00#, 16#00#, 16#10#, 16#00#, -- 33
		16#28#, 16#28#, 16#28#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, -- 34
		16#24#, 16#7e#, 16#24#, 16#24#, 16#24#, 16#7e#, 16#24#, 16#00#, -- 35
		16#10#, 16#3c#, 16#50#, 16#38#, 16#14#, 16#78#, 16#10#, 16#00#, -- 36
		16#60#, 16#64#, 16#08#, 16#10#, 16#20#, 16#4c#, 16#0c#, 16#00#, -- 37
		16#10#, 16#28#, 16#28#, 16#30#, 16#54#, 16#48#, 16#34#, 16#00#, -- 38
		16#10#, 16#10#, 16#20#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, -- 39
		16#08#, 16#10#, 16#20#, 16#20#, 16#20#, 16#10#, 16#08#, 16#00#, -- 40
		16#20#, 16#10#, 16#08#, 16#08#, 16#08#, 16#10#, 16#20#, 16#00#, -- 41
		16#00#, 16#10#, 16#54#, 16#38#, 16#54#, 16#10#, 16#00#, 16#00#, -- 42
		16#00#, 16#10#, 16#10#, 16#7c#, 16#10#, 16#10#, 16#00#, 16#00#, -- 43
		16#00#, 16#00#, 16#00#, 16#00#, 16#10#, 16#10#, 16#20#, 16#00#, -- 44
		16#00#, 16#00#, 16#00#, 16#7c#, 16#00#, 16#00#, 16#00#, 16#00#, -- 45
		16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#30#, 16#30#, 16#00#, -- 46
		16#00#, 16#04#, 16#08#, 16#10#, 16#20#, 16#40#, 16#00#, 16#00#, -- 47
		16#38#, 16#44#, 16#4c#, 16#54#, 16#64#, 16#44#, 16#38#, 16#00#, -- 48
		16#10#, 16#30#, 16#10#, 16#10#, 16#10#, 16#10#, 16#38#, 16#00#, -- 49
		16#38#, 16#44#, 16#04#, 16#08#, 16#10#, 16#20#, 16#7c#, 16#00#, -- 50
		16#7c#, 16#08#, 16#10#, 16#08#, 16#04#, 16#44#, 16#38#, 16#00#, -- 51
		16#08#, 16#18#, 16#28#, 16#48#, 16#7c#, 16#08#, 16#08#, 16#00#, -- 52
		16#7c#, 16#40#, 16#78#, 16#04#, 16#04#, 16#44#, 16#38#, 16#00#, -- 53
		16#18#, 16#20#, 16#40#, 16#78#, 16#44#, 16#44#, 16#38#, 16#00#, -- 54
		16#7c#, 16#04#, 16#08#, 16#10#, 16#20#, 16#20#, 16#20#, 16#00#, -- 55
		16#38#, 16#44#, 16#44#, 16#38#, 16#44#, 16#44#, 16#38#, 16#00#, -- 56
		16#38#, 16#44#, 16#44#, 16#3c#, 16#04#, 16#08#, 16#30#, 16#00#, -- 57
		16#00#, 16#30#, 16#30#, 16#00#, 16#30#, 16#30#, 16#00#, 16#00#, -- 58
		16#00#, 16#00#, 16#10#, 16#00#, 16#10#, 16#10#, 16#20#, 16#00#, -- 59
		16#08#, 16#10#, 16#20#, 16#40#, 16#20#, 16#10#, 16#08#, 16#00#, -- 60
		16#00#, 16#00#, 16#7c#, 16#00#, 16#7c#, 16#00#, 16#00#, 16#00#, -- 61
		16#20#, 16#10#, 16#08#, 16#04#, 16#08#, 16#10#, 16#20#, 16#00#, -- 62
		16#38#, 16#44#, 16#04#, 16#08#, 16#10#, 16#00#, 16#10#, 16#00#, -- 63
		16#38#, 16#44#, 16#5c#, 16#54#, 16#5c#, 16#40#, 16#3c#, 16#00#, -- 64
		16#38#, 16#44#, 16#44#, 16#7c#, 16#44#, 16#44#, 16#44#, 16#00#, -- 65
		16#78#, 16#24#, 16#24#, 16#38#, 16#24#, 16#24#, 16#78#, 16#00#, -- 66
		16#38#, 16#44#, 16#40#, 16#40#, 16#40#, 16#44#, 16#38#, 16#00#, -- 67
		16#78#, 16#24#, 16#24#, 16#24#, 16#24#, 16#24#, 16#78#, 16#00#, -- 68
		16#7c#, 16#40#, 16#40#, 16#78#, 16#40#, 16#40#, 16#7c#, 16#00#, -- 69
		16#7c#, 16#40#, 16#40#, 16#78#, 16#40#, 16#40#, 16#40#, 16#00#, -- 70
		16#38#, 16#44#, 16#40#, 16#40#, 16#4c#, 16#44#, 16#3c#, 16#00#, -- 71
		16#44#, 16#44#, 16#44#, 16#7c#, 16#44#, 16#44#, 16#44#, 16#00#, -- 72
		16#38#, 16#10#, 16#10#, 16#10#, 16#10#, 16#10#, 16#38#, 16#00#, -- 73
		16#1c#, 16#08#, 16#08#, 16#08#, 16#08#, 16#48#, 16#30#, 16#00#, -- 74
		16#44#, 16#48#, 16#50#, 16#60#, 16#50#, 16#48#, 16#44#, 16#00#, -- 75
		16#40#, 16#40#, 16#40#, 16#40#, 16#40#, 16#40#, 16#7c#, 16#00#, -- 76
		16#44#, 16#6c#, 16#54#, 16#54#, 16#44#, 16#44#, 16#44#, 16#00#, -- 77
		16#44#, 16#44#, 16#64#, 16#54#, 16#4c#, 16#44#, 16#44#, 16#00#, -- 78
		16#38#, 16#44#, 16#44#, 16#44#, 16#44#, 16#44#, 16#38#, 16#00#, -- 79
		16#78#, 16#44#, 16#44#, 16#78#, 16#40#, 16#40#, 16#40#, 16#00#, -- 80
		16#38#, 16#44#, 16#44#, 16#44#, 16#54#, 16#48#, 16#34#, 16#00#, -- 81
		16#78#, 16#44#, 16#44#, 16#78#, 16#50#, 16#48#, 16#44#, 16#00#, -- 82
		16#3c#, 16#40#, 16#40#, 16#38#, 16#04#, 16#04#, 16#78#, 16#00#, -- 83
		16#7c#, 16#10#, 16#10#, 16#10#, 16#10#, 16#10#, 16#10#, 16#00#, -- 84
		16#44#, 16#44#, 16#44#, 16#44#, 16#44#, 16#44#, 16#38#, 16#00#, -- 85
		16#44#, 16#44#, 16#44#, 16#44#, 16#44#, 16#28#, 16#10#, 16#00#, -- 86
		16#44#, 16#44#, 16#44#, 16#54#, 16#54#, 16#6c#, 16#44#, 16#00#, -- 87
		16#44#, 16#44#, 16#28#, 16#10#, 16#28#, 16#44#, 16#44#, 16#00#, -- 88
		16#44#, 16#44#, 16#44#, 16#28#, 16#10#, 16#10#, 16#10#, 16#00#, -- 89
		16#7c#, 16#04#, 16#08#, 16#10#, 16#20#, 16#40#, 16#7c#, 16#00#, -- 90
		16#44#, 16#38#, 16#44#, 16#44#, 16#7c#, 16#44#, 16#44#, 16#00#, -- 91
		16#44#, 16#38#, 16#44#, 16#44#, 16#44#, 16#44#, 16#38#, 16#00#, -- 92
		16#44#, 16#00#, 16#44#, 16#44#, 16#44#, 16#44#, 16#38#, 16#00#, -- 93
		16#10#, 16#28#, 16#44#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, -- 94
		16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#7e#, 16#00#, -- 95
		16#00#, 16#20#, 16#10#, 16#08#, 16#00#, 16#00#, 16#00#, 16#00#, -- 96
		16#00#, 16#00#, 16#34#, 16#4c#, 16#44#, 16#44#, 16#3a#, 16#00#, -- 97
		16#40#, 16#40#, 16#58#, 16#64#, 16#44#, 16#44#, 16#78#, 16#00#, -- 98
		16#00#, 16#00#, 16#38#, 16#44#, 16#40#, 16#44#, 16#38#, 16#00#, -- 99
		16#04#, 16#04#, 16#34#, 16#4c#, 16#44#, 16#44#, 16#3a#, 16#00#, -- 100
		16#00#, 16#00#, 16#38#, 16#44#, 16#7c#, 16#40#, 16#38#, 16#00#, -- 101
		16#08#, 16#10#, 16#38#, 16#10#, 16#10#, 16#10#, 16#10#, 16#00#, -- 102
		16#00#, 16#00#, 16#34#, 16#4c#, 16#44#, 16#3c#, 16#04#, 16#38#, -- 103
		16#40#, 16#40#, 16#58#, 16#64#, 16#44#, 16#44#, 16#44#, 16#00#, -- 104
		16#10#, 16#00#, 16#10#, 16#10#, 16#10#, 16#10#, 16#08#, 16#00#, -- 105
		16#10#, 16#00#, 16#10#, 16#10#, 16#10#, 16#10#, 16#10#, 16#20#, -- 106
		16#40#, 16#40#, 16#48#, 16#50#, 16#70#, 16#48#, 16#44#, 16#00#, -- 107
		16#10#, 16#10#, 16#10#, 16#10#, 16#10#, 16#10#, 16#08#, 16#00#, -- 108
		16#00#, 16#00#, 16#68#, 16#54#, 16#54#, 16#54#, 16#54#, 16#00#, -- 109
		16#00#, 16#00#, 16#58#, 16#64#, 16#44#, 16#44#, 16#44#, 16#00#, -- 110
		16#00#, 16#00#, 16#38#, 16#44#, 16#44#, 16#44#, 16#38#, 16#00#, -- 111
		16#00#, 16#00#, 16#58#, 16#64#, 16#44#, 16#78#, 16#40#, 16#40#, -- 112
		16#00#, 16#00#, 16#34#, 16#4c#, 16#44#, 16#3c#, 16#04#, 16#04#, -- 113
		16#00#, 16#00#, 16#58#, 16#64#, 16#40#, 16#40#, 16#40#, 16#00#, -- 114
		16#00#, 16#00#, 16#38#, 16#40#, 16#38#, 16#04#, 16#78#, 16#00#, -- 115
		16#10#, 16#10#, 16#38#, 16#10#, 16#10#, 16#10#, 16#08#, 16#00#, -- 116
		16#00#, 16#00#, 16#44#, 16#44#, 16#44#, 16#4c#, 16#34#, 16#00#, -- 117
		16#00#, 16#00#, 16#44#, 16#44#, 16#44#, 16#28#, 16#10#, 16#00#, -- 118
		16#00#, 16#00#, 16#54#, 16#54#, 16#54#, 16#54#, 16#28#, 16#00#, -- 119
		16#00#, 16#00#, 16#44#, 16#28#, 16#10#, 16#28#, 16#44#, 16#00#, -- 120
		16#00#, 16#00#, 16#44#, 16#44#, 16#44#, 16#3c#, 16#04#, 16#38#, -- 121
		16#00#, 16#00#, 16#7c#, 16#08#, 16#10#, 16#20#, 16#7c#, 16#00#, -- 122
		16#28#, 16#00#, 16#34#, 16#4c#, 16#44#, 16#44#, 16#3a#, 16#00#, -- 123
		16#28#, 16#00#, 16#38#, 16#44#, 16#44#, 16#44#, 16#38#, 16#00#, -- 124
		16#28#, 16#00#, 16#44#, 16#44#, 16#44#, 16#4c#, 16#34#, 16#00#, -- 125
		16#18#, 16#24#, 16#24#, 16#28#, 16#24#, 16#34#, 16#28#, 16#00#, -- 126
		16#ff#, 16#cf#, 16#e7#, 16#f3#, 16#e7#, 16#cf#, 16#ff#, 16#00#, -- 127
		16#ff#, 16#bb#, 16#55#, 16#55#, 16#55#, 16#55#, 16#bb#, 16#ff#, -- 128
		16#bf#, 16#5f#, 16#f3#, 16#ed#, 16#e1#, 16#ed#, 16#ed#, 16#ff#, -- 129
		16#bf#, 16#5f#, 16#e3#, 16#ed#, 16#e3#, 16#ed#, 16#e3#, 16#ff#, -- 130
		16#bf#, 16#5f#, 16#f3#, 16#ed#, 16#ef#, 16#ed#, 16#f3#, 16#ff#, -- 131
		16#bf#, 16#5f#, 16#e3#, 16#ed#, 16#ed#, 16#ed#, 16#e3#, 16#ff#, -- 132
		16#bf#, 16#5f#, 16#e1#, 16#ef#, 16#e3#, 16#ef#, 16#e1#, 16#ff#, -- 133
		16#bf#, 16#5f#, 16#e1#, 16#ef#, 16#e3#, 16#ef#, 16#ef#, 16#ff#, -- 134
		16#bf#, 16#5f#, 16#f3#, 16#ed#, 16#ef#, 16#e9#, 16#f1#, 16#ff#, -- 135
		16#bf#, 16#5f#, 16#ed#, 16#ed#, 16#e1#, 16#ed#, 16#ed#, 16#ff#, -- 136
		16#bf#, 16#5f#, 16#f1#, 16#fb#, 16#fb#, 16#fb#, 16#f1#, 16#ff#, -- 137
		16#ff#, 16#ff#, 16#71#, 16#77#, 16#73#, 16#77#, 16#17#, 16#ff#, -- 138
		16#bf#, 16#5f#, 16#ed#, 16#eb#, 16#e7#, 16#eb#, 16#ed#, 16#ff#, -- 139
		16#bf#, 16#5f#, 16#ef#, 16#ef#, 16#ef#, 16#ef#, 16#e1#, 16#ff#, -- 140
		16#ff#, 16#ff#, 16#93#, 16#75#, 16#73#, 16#75#, 16#95#, 16#ff#, -- 141
		16#bf#, 16#5f#, 16#ed#, 16#e5#, 16#e9#, 16#ed#, 16#ed#, 16#ff#, -- 142
		16#bf#, 16#5f#, 16#f3#, 16#ed#, 16#ed#, 16#ed#, 16#f3#, 16#ff#, -- 143
		16#bf#, 16#5f#, 16#e3#, 16#ed#, 16#e3#, 16#ef#, 16#ef#, 16#ff#, -- 144
		16#bf#, 16#5f#, 16#f3#, 16#ed#, 16#ed#, 16#eb#, 16#f5#, 16#ff#, -- 145
		16#bf#, 16#5f#, 16#e3#, 16#ed#, 16#e3#, 16#eb#, 16#ed#, 16#ff#, -- 146
		16#bf#, 16#5f#, 16#f1#, 16#ef#, 16#f3#, 16#fd#, 16#e3#, 16#ff#, -- 147
		16#bf#, 16#5f#, 16#f1#, 16#fb#, 16#fb#, 16#fb#, 16#fb#, 16#ff#, -- 148
		16#bf#, 16#5f#, 16#ed#, 16#ed#, 16#ed#, 16#ed#, 16#f3#, 16#ff#, -- 149
		16#bf#, 16#5f#, 16#ee#, 16#ee#, 16#ee#, 16#f5#, 16#fb#, 16#ff#, -- 150
		16#bf#, 16#5f#, 16#ee#, 16#ea#, 16#ea#, 16#e4#, 16#ee#, 16#ff#, -- 151
		16#bf#, 16#5f#, 16#ee#, 16#f5#, 16#fb#, 16#f5#, 16#ee#, 16#ff#, -- 152
		16#bf#, 16#5f#, 16#ee#, 16#ee#, 16#f5#, 16#fb#, 16#fb#, 16#ff#, -- 153
		16#bf#, 16#5f#, 16#e1#, 16#fd#, 16#fb#, 16#f7#, 16#e1#, 16#ff#, -- 154
		16#ff#, 16#ff#, 16#24#, 16#6d#, 16#35#, 16#75#, 16#24#, 16#ff#, -- 155
		16#b7#, 16#57#, 16#f7#, 16#f7#, 16#f7#, 16#f7#, 16#ff#, 16#ff#, -- 156
		16#bf#, 16#5f#, 16#f3#, 16#fb#, 16#f9#, 16#fb#, 16#f3#, 16#ff#, -- 157
		16#ff#, 16#ff#, 16#6b#, 16#2b#, 16#4b#, 16#6b#, 16#69#, 16#ff#, -- 158
		16#ff#, 16#ff#, 16#d1#, 16#97#, 16#d3#, 16#d7#, 16#d7#, 16#ff#, -- 159
		16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, -- 160
		16#ef#, 16#ef#, 16#ef#, 16#ef#, 16#ff#, 16#ff#, 16#ef#, 16#ff#, -- 161
		16#d7#, 16#d7#, 16#d7#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, -- 162
		16#db#, 16#81#, 16#db#, 16#db#, 16#db#, 16#81#, 16#db#, 16#ff#, -- 163
		16#ef#, 16#c3#, 16#af#, 16#c7#, 16#eb#, 16#87#, 16#ef#, 16#ff#, -- 164
		16#9f#, 16#9b#, 16#f7#, 16#ef#, 16#df#, 16#b3#, 16#f3#, 16#ff#, -- 165
		16#ef#, 16#d7#, 16#d7#, 16#cf#, 16#ab#, 16#b7#, 16#cb#, 16#ff#, -- 166
		16#ef#, 16#ef#, 16#df#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, -- 167
		16#f7#, 16#ef#, 16#df#, 16#df#, 16#df#, 16#ef#, 16#f7#, 16#ff#, -- 168
		16#df#, 16#ef#, 16#f7#, 16#f7#, 16#f7#, 16#ef#, 16#df#, 16#ff#, -- 169
		16#ff#, 16#ef#, 16#ab#, 16#c7#, 16#ab#, 16#ef#, 16#ff#, 16#ff#, -- 170
		16#ff#, 16#ef#, 16#ef#, 16#83#, 16#ef#, 16#ef#, 16#ff#, 16#ff#, -- 171
		16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ef#, 16#ef#, 16#df#, 16#ff#, -- 172
		16#ff#, 16#ff#, 16#ff#, 16#83#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, -- 173
		16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#cf#, 16#cf#, 16#ff#, -- 174
		16#ff#, 16#fb#, 16#f7#, 16#ef#, 16#df#, 16#bf#, 16#ff#, 16#ff#, -- 175
		16#c7#, 16#bb#, 16#b3#, 16#ab#, 16#9b#, 16#bb#, 16#c7#, 16#ff#, -- 176
		16#ef#, 16#cf#, 16#ef#, 16#ef#, 16#ef#, 16#ef#, 16#c7#, 16#ff#, -- 177
		16#c7#, 16#bb#, 16#fb#, 16#f7#, 16#ef#, 16#df#, 16#83#, 16#ff#, -- 178
		16#83#, 16#f7#, 16#ef#, 16#f7#, 16#fb#, 16#bb#, 16#c7#, 16#ff#, -- 179
		16#f7#, 16#e7#, 16#d7#, 16#b7#, 16#83#, 16#f7#, 16#f7#, 16#ff#, -- 180
		16#83#, 16#bf#, 16#87#, 16#fb#, 16#fb#, 16#bb#, 16#c7#, 16#ff#, -- 181
		16#e7#, 16#df#, 16#bf#, 16#87#, 16#bb#, 16#bb#, 16#c7#, 16#ff#, -- 182
		16#83#, 16#fb#, 16#f7#, 16#ef#, 16#df#, 16#df#, 16#df#, 16#ff#, -- 183
		16#c7#, 16#bb#, 16#bb#, 16#c7#, 16#bb#, 16#bb#, 16#c7#, 16#ff#, -- 184
		16#c7#, 16#bb#, 16#bb#, 16#c3#, 16#fb#, 16#f7#, 16#cf#, 16#ff#, -- 185
		16#ff#, 16#cf#, 16#cf#, 16#ff#, 16#cf#, 16#cf#, 16#ff#, 16#ff#, -- 186
		16#ff#, 16#ff#, 16#ef#, 16#ff#, 16#ef#, 16#ef#, 16#df#, 16#ff#, -- 187
		16#f7#, 16#ef#, 16#df#, 16#bf#, 16#df#, 16#ef#, 16#f7#, 16#ff#, -- 188
		16#ff#, 16#ff#, 16#83#, 16#ff#, 16#83#, 16#ff#, 16#ff#, 16#ff#, -- 189
		16#df#, 16#ef#, 16#f7#, 16#fb#, 16#f7#, 16#ef#, 16#df#, 16#ff#, -- 190
		16#c7#, 16#bb#, 16#fb#, 16#f7#, 16#ef#, 16#ff#, 16#ef#, 16#ff#, -- 191
		16#c7#, 16#bb#, 16#a3#, 16#ab#, 16#a3#, 16#bf#, 16#c3#, 16#ff#, -- 192
		16#c7#, 16#bb#, 16#bb#, 16#83#, 16#bb#, 16#bb#, 16#bb#, 16#ff#, -- 193
		16#87#, 16#db#, 16#db#, 16#c7#, 16#db#, 16#db#, 16#87#, 16#ff#, -- 194
		16#c7#, 16#bb#, 16#bf#, 16#bf#, 16#bf#, 16#bb#, 16#c7#, 16#ff#, -- 195
		16#87#, 16#db#, 16#db#, 16#db#, 16#db#, 16#db#, 16#87#, 16#ff#, -- 196
		16#83#, 16#bf#, 16#bf#, 16#87#, 16#bf#, 16#bf#, 16#83#, 16#ff#, -- 197
		16#83#, 16#bf#, 16#bf#, 16#87#, 16#bf#, 16#bf#, 16#bf#, 16#ff#, -- 198
		16#c7#, 16#bb#, 16#bf#, 16#bf#, 16#b3#, 16#bb#, 16#c3#, 16#ff#, -- 199
		16#bb#, 16#bb#, 16#bb#, 16#83#, 16#bb#, 16#bb#, 16#bb#, 16#ff#, -- 200
		16#c7#, 16#ef#, 16#ef#, 16#ef#, 16#ef#, 16#ef#, 16#c7#, 16#ff#, -- 201
		16#e3#, 16#f7#, 16#f7#, 16#f7#, 16#f7#, 16#b7#, 16#cf#, 16#ff#, -- 202
		16#bb#, 16#b7#, 16#af#, 16#9f#, 16#af#, 16#b7#, 16#bb#, 16#ff#, -- 203
		16#bf#, 16#bf#, 16#bf#, 16#bf#, 16#bf#, 16#bf#, 16#83#, 16#ff#, -- 204
		16#bb#, 16#93#, 16#ab#, 16#ab#, 16#bb#, 16#bb#, 16#bb#, 16#ff#, -- 205
		16#bb#, 16#bb#, 16#9b#, 16#ab#, 16#b3#, 16#bb#, 16#bb#, 16#ff#, -- 206
		16#c7#, 16#bb#, 16#bb#, 16#bb#, 16#bb#, 16#bb#, 16#c7#, 16#ff#, -- 207
		16#87#, 16#bb#, 16#bb#, 16#87#, 16#bf#, 16#bf#, 16#bf#, 16#ff#, -- 208
		16#c7#, 16#bb#, 16#bb#, 16#bb#, 16#ab#, 16#b7#, 16#cb#, 16#ff#, -- 209
		16#87#, 16#bb#, 16#bb#, 16#87#, 16#af#, 16#b7#, 16#bb#, 16#ff#, -- 210
		16#c3#, 16#bf#, 16#bf#, 16#c7#, 16#fb#, 16#fb#, 16#87#, 16#ff#, -- 211
		16#83#, 16#ef#, 16#ef#, 16#ef#, 16#ef#, 16#ef#, 16#ef#, 16#ff#, -- 212
		16#bb#, 16#bb#, 16#bb#, 16#bb#, 16#bb#, 16#bb#, 16#c7#, 16#ff#, -- 213
		16#bb#, 16#bb#, 16#bb#, 16#bb#, 16#bb#, 16#d7#, 16#ef#, 16#ff#, -- 214
		16#bb#, 16#bb#, 16#bb#, 16#ab#, 16#ab#, 16#93#, 16#bb#, 16#ff#, -- 215
		16#bb#, 16#bb#, 16#d7#, 16#ef#, 16#d7#, 16#bb#, 16#bb#, 16#ff#, -- 216
		16#bb#, 16#bb#, 16#bb#, 16#d7#, 16#ef#, 16#ef#, 16#ef#, 16#ff#, -- 217
		16#83#, 16#fb#, 16#f7#, 16#ef#, 16#df#, 16#bf#, 16#83#, 16#ff#, -- 218
		16#bb#, 16#c7#, 16#bb#, 16#bb#, 16#83#, 16#bb#, 16#bb#, 16#ff#, -- 219
		16#bb#, 16#c7#, 16#bb#, 16#bb#, 16#bb#, 16#bb#, 16#c7#, 16#ff#, -- 220
		16#bb#, 16#ff#, 16#bb#, 16#bb#, 16#bb#, 16#bb#, 16#c7#, 16#ff#, -- 221
		16#ef#, 16#d7#, 16#bb#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, -- 222
		16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#81#, 16#ff#, -- 223
		16#ff#, 16#df#, 16#ef#, 16#f7#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, -- 224
		16#ff#, 16#ff#, 16#cb#, 16#b3#, 16#bb#, 16#bb#, 16#c5#, 16#ff#, -- 225
		16#bf#, 16#bf#, 16#a7#, 16#9b#, 16#bb#, 16#bb#, 16#87#, 16#ff#, -- 226
		16#ff#, 16#ff#, 16#c7#, 16#bb#, 16#bf#, 16#bb#, 16#c7#, 16#ff#, -- 227
		16#fb#, 16#fb#, 16#cb#, 16#b3#, 16#bb#, 16#bb#, 16#c5#, 16#ff#, -- 228
		16#ff#, 16#ff#, 16#c7#, 16#bb#, 16#83#, 16#bf#, 16#c7#, 16#ff#, -- 229
		16#f7#, 16#ef#, 16#c7#, 16#ef#, 16#ef#, 16#ef#, 16#ef#, 16#ff#, -- 230
		16#ff#, 16#ff#, 16#cb#, 16#b3#, 16#bb#, 16#c3#, 16#fb#, 16#c7#, -- 231
		16#bf#, 16#bf#, 16#a7#, 16#9b#, 16#bb#, 16#bb#, 16#bb#, 16#ff#, -- 232
		16#ef#, 16#ff#, 16#ef#, 16#ef#, 16#ef#, 16#ef#, 16#f7#, 16#ff#, -- 233
		16#ef#, 16#ff#, 16#ef#, 16#ef#, 16#ef#, 16#ef#, 16#ef#, 16#df#, -- 234
		16#bf#, 16#bf#, 16#b7#, 16#af#, 16#8f#, 16#b7#, 16#bb#, 16#ff#, -- 235
		16#ef#, 16#ef#, 16#ef#, 16#ef#, 16#ef#, 16#ef#, 16#f7#, 16#ff#, -- 236
		16#ff#, 16#ff#, 16#97#, 16#ab#, 16#ab#, 16#ab#, 16#ab#, 16#ff#, -- 237
		16#ff#, 16#ff#, 16#a7#, 16#9b#, 16#bb#, 16#bb#, 16#bb#, 16#ff#, -- 238
		16#ff#, 16#ff#, 16#c7#, 16#bb#, 16#bb#, 16#bb#, 16#c7#, 16#ff#, -- 239
		16#ff#, 16#ff#, 16#a7#, 16#9b#, 16#bb#, 16#87#, 16#bf#, 16#bf#, -- 240
		16#ff#, 16#ff#, 16#cb#, 16#b3#, 16#bb#, 16#c3#, 16#fb#, 16#fb#, -- 241
		16#ff#, 16#ff#, 16#a7#, 16#9b#, 16#bf#, 16#bf#, 16#bf#, 16#ff#, -- 242
		16#ff#, 16#ff#, 16#c7#, 16#bf#, 16#c7#, 16#fb#, 16#87#, 16#ff#, -- 243
		16#ef#, 16#ef#, 16#c7#, 16#ef#, 16#ef#, 16#ef#, 16#f7#, 16#ff#, -- 244
		16#ff#, 16#ff#, 16#bb#, 16#bb#, 16#bb#, 16#b3#, 16#cb#, 16#ff#, -- 245
		16#ff#, 16#ff#, 16#bb#, 16#bb#, 16#bb#, 16#d7#, 16#ef#, 16#ff#, -- 246
		16#ff#, 16#ff#, 16#ab#, 16#ab#, 16#ab#, 16#ab#, 16#d7#, 16#ff#, -- 247
		16#ff#, 16#ff#, 16#bb#, 16#d7#, 16#ef#, 16#d7#, 16#bb#, 16#ff#, -- 248
		16#ff#, 16#ff#, 16#bb#, 16#bb#, 16#bb#, 16#c3#, 16#fb#, 16#c7#, -- 249
		16#ff#, 16#ff#, 16#83#, 16#f7#, 16#ef#, 16#df#, 16#83#, 16#ff#, -- 250
		16#d7#, 16#ff#, 16#cb#, 16#b3#, 16#bb#, 16#bb#, 16#c5#, 16#ff#, -- 251
		16#d7#, 16#ff#, 16#c7#, 16#bb#, 16#bb#, 16#bb#, 16#c7#, 16#ff#, -- 252
		16#d7#, 16#ff#, 16#bb#, 16#bb#, 16#bb#, 16#b3#, 16#cb#, 16#ff#, -- 253
		16#e7#, 16#db#, 16#db#, 16#d7#, 16#db#, 16#cb#, 16#d7#, 16#ff#, -- 254
		16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#  -- 255
    );

    signal crom_array : T_BM100_MEM := charrom2_init;
    signal crom_index : natural;


begin

    crom_index <= to_integer( unsigned( addr_char_i & addr_line_i));
  
    process
    begin
        wait until rising_edge( clk);
        data_o <= std_logic_vector( to_unsigned( crom_array( crom_index), 8));
    end process;

end architecture rtl;
