------------------------------------------------------------------------------
-- Project    : Red Zombie
------------------------------------------------------------------------------
-- File       :  bm100_pkg.vhd
-- Author     :  fpgakuechle
-- Company    : hobbyist
-- Created    : 2012-12
-- Last update: 2013-06-30
-- Licence    : 
------------------------------------------------------------------------------
-- Description: 
-- converted rom image
-- Z1013 EPROM-image U2632  bm100 Bitmuster 100
-- char set (numbers,letters, graphic symbols, chess figures, .. 
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

package bm100_pkg is
  subtype T_BM100_INDEX is integer range 0 to 2**11 - 1;
  subtype T_WORD is integer range 255 downto 0;
  type    T_BM100_MEM is array (T_BM100_INDEX'low to T_BM100_INDEX'high) of T_word;

--'0' - '9' x30 -x39
--'A' - 'F' x41 -x46  
--'a' - 'f' x61 -x66  
constant C_BM100_MEM_ARRAY_INIT : T_BM100_MEM := (
16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#,--x00|x01
16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#,
16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#,
16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#,
16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#,--x08|x09
16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#,
16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#,--x0c|0D
16#00#, 16#00#, 16#18#, 16#24#, 16#24#, 16#18#, 16#24#, 16#42#, 16#db#, 16#a5#, 16#81#, 16#ff#, 16#24#, 16#24#, 16#24#, 16#42#,--x0E|x0F chess piece 
16#08#, 16#34#, 16#42#, 16#81#, 16#91#, 16#69#, 16#09#, 16#31#, 16#42#, 16#7e#, 16#81#, 16#ff#, 16#00#, 16#00#, 16#00#, 16#00#,  --x10
16#18#, 16#24#, 16#42#, 16#99#, 16#bd#, 16#99#, 16#42#, 16#24#, 16#7e#, 16#42#, 16#99#, 16#e7#, 16#00#, 16#00#, 16#00#, 16#00#,
16#18#, 16#db#, 16#c3#, 16#18#, 16#99#, 16#e7#, 16#81#, 16#42#, 16#18#, 16#24#, 16#18#, 16#c3#, 16#bd#, 16#81#, 16#81#, 16#42#,
16#24#, 16#7e#, 16#81#, 16#ff#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#18#, 16#3c#, 16#3c#, 16#18#, 16#3c#, 16#7e#,
16#db#, 16#ff#, 16#ff#, 16#ff#, 16#3c#, 16#3c#, 16#3c#, 16#7e#, 16#08#, 16#3c#, 16#7e#, 16#ff#, 16#ff#, 16#6f#, 16#0f#, 16#3f#, -- x18
16#7e#, 16#7e#, 16#ff#, 16#ff#, 16#00#, 16#00#, 16#00#, 16#00#, 16#18#, 16#3c#, 16#7e#, 16#e7#, 16#c3#, 16#e7#, 16#7e#, 16#3c#,
16#7e#, 16#7e#, 16#ff#, 16#e7#, 16#00#, 16#00#, 16#00#, 16#00#, 16#18#, 16#db#, 16#c3#, 16#18#, 16#99#, 16#ff#, 16#ff#, 16#7e#,
16#18#, 16#3c#, 16#18#, 16#c3#, 16#ff#, 16#ff#, 16#ff#, 16#7e#, 16#3c#, 16#3c#, 16#ff#, 16#ff#, 16#00#, 16#00#, 16#00#, 16#00#,
16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#10#, 16#10#, 16#10#, 16#10#, 16#00#, 16#00#, 16#10#, 16#00#,--x20|x21 space+'!'
16#28#, 16#28#, 16#28#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#24#, 16#7e#, 16#24#, 16#24#, 16#24#, 16#7e#, 16#24#, 16#00#,
16#10#, 16#3c#, 16#50#, 16#38#, 16#14#, 16#78#, 16#10#, 16#00#, 16#60#, 16#64#, 16#08#, 16#10#, 16#20#, 16#4c#, 16#0c#, 16#00#,
16#10#, 16#28#, 16#28#, 16#30#, 16#54#, 16#48#, 16#34#, 16#00#, 16#10#, 16#10#, 16#20#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#,
16#08#, 16#10#, 16#20#, 16#20#, 16#20#, 16#10#, 16#08#, 16#00#, 16#20#, 16#10#, 16#08#, 16#08#, 16#08#, 16#10#, 16#20#, 16#00#, -- x28
16#00#, 16#10#, 16#54#, 16#38#, 16#54#, 16#10#, 16#00#, 16#00#, 16#00#, 16#10#, 16#10#, 16#7c#, 16#10#, 16#10#, 16#00#, 16#00#,
16#00#, 16#00#, 16#00#, 16#00#, 16#10#, 16#10#, 16#20#, 16#00#, 16#00#, 16#00#, 16#00#, 16#7c#, 16#00#, 16#00#, 16#00#, 16#00#,
16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#30#, 16#30#, 16#00#, 16#00#, 16#04#, 16#08#, 16#10#, 16#20#, 16#40#, 16#00#, 16#00#,
16#38#, 16#44#, 16#44#, 16#54#, 16#44#, 16#44#, 16#38#, 16#00#, 16#10#, 16#30#, 16#10#, 16#10#, 16#10#, 16#10#, 16#38#, 16#00#,--x30 0 1
16#38#, 16#44#, 16#04#, 16#08#, 16#10#, 16#20#, 16#7c#, 16#00#, 16#7c#, 16#08#, 16#10#, 16#08#, 16#04#, 16#44#, 16#38#, 16#00#,--2 3
16#08#, 16#18#, 16#28#, 16#48#, 16#7c#, 16#08#, 16#08#, 16#00#, 16#7c#, 16#40#, 16#78#, 16#04#, 16#04#, 16#44#, 16#38#, 16#00#,-- 4 5
16#18#, 16#20#, 16#40#, 16#78#, 16#44#, 16#44#, 16#38#, 16#00#, 16#7c#, 16#04#, 16#08#, 16#10#, 16#20#, 16#20#, 16#20#, 16#00#,-- 6 7
16#38#, 16#44#, 16#44#, 16#38#, 16#44#, 16#44#, 16#38#, 16#00#, 16#38#, 16#44#, 16#44#, 16#3c#, 16#04#, 16#08#, 16#30#, 16#00#,-- 8 9
16#00#, 16#30#, 16#30#, 16#00#, 16#30#, 16#30#, 16#00#, 16#00#, 16#00#, 16#00#, 16#10#, 16#00#, 16#10#, 16#10#, 16#20#, 16#00#,
16#08#, 16#10#, 16#20#, 16#40#, 16#20#, 16#10#, 16#08#, 16#00#, 16#00#, 16#00#, 16#7c#, 16#00#, 16#7c#, 16#00#, 16#00#, 16#00#,
16#20#, 16#10#, 16#08#, 16#04#, 16#08#, 16#10#, 16#20#, 16#00#, 16#38#, 16#44#, 16#04#, 16#08#, 16#10#, 16#00#, 16#10#, 16#00#,
16#38#, 16#44#, 16#5c#, 16#54#, 16#5c#, 16#40#, 16#3c#, 16#00#, 16#38#, 16#44#, 16#44#, 16#7c#, 16#44#, 16#44#, 16#44#, 16#00#,--x40 @ A
16#78#, 16#24#, 16#24#, 16#38#, 16#24#, 16#24#, 16#78#, 16#00#, 16#38#, 16#44#, 16#40#, 16#40#, 16#40#, 16#44#, 16#38#, 16#00#,-- B C
16#78#, 16#24#, 16#24#, 16#24#, 16#24#, 16#24#, 16#78#, 16#00#, 16#7c#, 16#40#, 16#40#, 16#78#, 16#40#, 16#40#, 16#7c#, 16#00#,-- D E
16#7c#, 16#40#, 16#40#, 16#78#, 16#40#, 16#40#, 16#40#, 16#00#, 16#38#, 16#44#, 16#40#, 16#40#, 16#4c#, 16#44#, 16#3c#, 16#00#,-- F G
16#44#, 16#44#, 16#44#, 16#7c#, 16#44#, 16#44#, 16#44#, 16#00#, 16#38#, 16#10#, 16#10#, 16#10#, 16#10#, 16#10#, 16#38#, 16#00#, -- x48
16#1c#, 16#08#, 16#08#, 16#08#, 16#08#, 16#48#, 16#30#, 16#00#, 16#44#, 16#48#, 16#50#, 16#60#, 16#50#, 16#48#, 16#44#, 16#00#,
16#40#, 16#40#, 16#40#, 16#40#, 16#40#, 16#40#, 16#7c#, 16#00#, 16#44#, 16#6c#, 16#54#, 16#54#, 16#44#, 16#44#, 16#44#, 16#00#,
16#44#, 16#44#, 16#64#, 16#54#, 16#4c#, 16#44#, 16#44#, 16#00#, 16#38#, 16#44#, 16#44#, 16#44#, 16#44#, 16#44#, 16#38#, 16#00#,
16#78#, 16#44#, 16#44#, 16#78#, 16#40#, 16#40#, 16#40#, 16#00#, 16#38#, 16#44#, 16#44#, 16#44#, 16#54#, 16#48#, 16#34#, 16#00#,--x50
16#78#, 16#44#, 16#44#, 16#78#, 16#50#, 16#48#, 16#44#, 16#00#, 16#3c#, 16#40#, 16#40#, 16#38#, 16#04#, 16#04#, 16#78#, 16#00#,
16#7c#, 16#10#, 16#10#, 16#10#, 16#10#, 16#10#, 16#10#, 16#00#, 16#44#, 16#44#, 16#44#, 16#44#, 16#44#, 16#44#, 16#38#, 16#00#,
16#44#, 16#44#, 16#44#, 16#44#, 16#44#, 16#28#, 16#10#, 16#00#, 16#44#, 16#44#, 16#44#, 16#54#, 16#54#, 16#6c#, 16#44#, 16#00#,
16#44#, 16#44#, 16#28#, 16#10#, 16#28#, 16#44#, 16#44#, 16#00#, 16#44#, 16#44#, 16#44#, 16#28#, 16#10#, 16#10#, 16#10#, 16#00#, -- x58
16#7c#, 16#04#, 16#08#, 16#10#, 16#20#, 16#40#, 16#7c#, 16#00#, 16#38#, 16#20#, 16#20#, 16#20#, 16#20#, 16#20#, 16#38#, 16#00#,
16#00#, 16#40#, 16#20#, 16#10#, 16#08#, 16#04#, 16#00#, 16#00#, 16#38#, 16#08#, 16#08#, 16#08#, 16#08#, 16#08#, 16#38#, 16#00#,
16#10#, 16#28#, 16#44#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#7c#, 16#00#, 16#00#,
16#00#, 16#20#, 16#10#, 16#08#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#34#, 16#4c#, 16#44#, 16#44#, 16#3a#, 16#00#, --x60 ' a 
16#40#, 16#40#, 16#58#, 16#64#, 16#44#, 16#44#, 16#78#, 16#00#, 16#00#, 16#00#, 16#38#, 16#44#, 16#40#, 16#44#, 16#38#, 16#00#, -- b c
16#04#, 16#04#, 16#34#, 16#4c#, 16#44#, 16#44#, 16#3a#, 16#00#, 16#00#, 16#00#, 16#38#, 16#44#, 16#7c#, 16#40#, 16#38#, 16#00#, -- d e
16#08#, 16#10#, 16#38#, 16#10#, 16#10#, 16#10#, 16#10#, 16#00#, 16#00#, 16#00#, 16#34#, 16#4c#, 16#44#, 16#3c#, 16#04#, 16#38#, -- f g
16#40#, 16#40#, 16#58#, 16#64#, 16#44#, 16#44#, 16#44#, 16#00#, 16#10#, 16#00#, 16#10#, 16#10#, 16#10#, 16#10#, 16#08#, 16#00#, -- x68
16#10#, 16#00#, 16#10#, 16#10#, 16#10#, 16#10#, 16#10#, 16#20#, 16#40#, 16#40#, 16#48#, 16#50#, 16#70#, 16#48#, 16#44#, 16#00#,
16#10#, 16#10#, 16#10#, 16#10#, 16#10#, 16#10#, 16#08#, 16#00#, 16#00#, 16#00#, 16#68#, 16#54#, 16#54#, 16#54#, 16#54#, 16#00#,
16#00#, 16#00#, 16#58#, 16#64#, 16#44#, 16#44#, 16#44#, 16#00#, 16#00#, 16#00#, 16#38#, 16#44#, 16#44#, 16#44#, 16#38#, 16#00#,
16#00#, 16#00#, 16#58#, 16#64#, 16#44#, 16#78#, 16#40#, 16#40#, 16#00#, 16#00#, 16#34#, 16#4c#, 16#44#, 16#3c#, 16#04#, 16#04#, -- x70
16#00#, 16#00#, 16#58#, 16#64#, 16#40#, 16#40#, 16#40#, 16#00#, 16#00#, 16#00#, 16#38#, 16#40#, 16#38#, 16#04#, 16#78#, 16#00#,
16#10#, 16#10#, 16#38#, 16#10#, 16#10#, 16#10#, 16#08#, 16#00#, 16#00#, 16#00#, 16#44#, 16#44#, 16#44#, 16#4c#, 16#34#, 16#00#,
16#00#, 16#00#, 16#44#, 16#44#, 16#44#, 16#28#, 16#10#, 16#00#, 16#00#, 16#00#, 16#54#, 16#54#, 16#54#, 16#54#, 16#28#, 16#00#,
16#00#, 16#00#, 16#44#, 16#28#, 16#10#, 16#28#, 16#44#, 16#00#, 16#00#, 16#00#, 16#44#, 16#44#, 16#44#, 16#3c#, 16#04#, 16#38#, -- x78
16#00#, 16#00#, 16#7c#, 16#08#, 16#10#, 16#20#, 16#7c#, 16#00#, 16#08#, 16#10#, 16#10#, 16#20#, 16#10#, 16#10#, 16#08#, 16#00#,
16#10#, 16#10#, 16#10#, 16#10#, 16#10#, 16#10#, 16#10#, 16#00#, 16#20#, 16#10#, 16#10#, 16#08#, 16#10#, 16#10#, 16#20#, 16#00#,
16#00#, 16#00#, 16#00#, 16#32#, 16#4c#, 16#00#, 16#00#, 16#00#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#,
16#c0#, 16#20#, 16#10#, 16#10#, 16#10#, 16#10#, 16#20#, 16#c0#, 16#03#, 16#04#, 16#08#, 16#08#, 16#08#, 16#08#, 16#04#, 16#03#, -- x80
16#81#, 16#81#, 16#42#, 16#3c#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#3c#, 16#42#, 16#81#, 16#81#,
16#10#, 16#10#, 16#20#, 16#c0#, 16#00#, 16#00#, 16#00#, 16#00#, 16#08#, 16#08#, 16#04#, 16#03#, 16#00#, 16#00#, 16#00#, 16#00#,
16#00#, 16#00#, 16#00#, 16#00#, 16#03#, 16#04#, 16#08#, 16#08#, 16#00#, 16#00#, 16#00#, 16#00#, 16#c0#, 16#20#, 16#10#, 16#10#,
16#80#, 16#80#, 16#80#, 16#80#, 16#80#, 16#80#, 16#80#, 16#ff#, 16#ff#, 16#01#, 16#01#, 16#01#, 16#01#, 16#01#, 16#01#, 16#01#, -- x88
16#00#, 16#10#, 16#28#, 16#44#, 16#82#, 16#44#, 16#28#, 16#10#, 16#ff#, 16#ef#, 16#c7#, 16#83#, 16#01#, 16#83#, 16#c7#, 16#ef#,
16#3c#, 16#42#, 16#81#, 16#81#, 16#81#, 16#81#, 16#42#, 16#3c#, 16#c3#, 16#81#, 16#00#, 16#00#, 16#00#, 16#00#, 16#81#, 16#c3#,
16#ff#, 16#fe#, 16#fc#, 16#f8#, 16#f0#, 16#e0#, 16#c0#, 16#80#, 16#80#, 16#c0#, 16#e0#, 16#f0#, 16#f8#, 16#fc#, 16#fe#, 16#ff#,
16#01#, 16#02#, 16#04#, 16#08#, 16#10#, 16#20#, 16#40#, 16#80#, 16#80#, 16#40#, 16#20#, 16#10#, 16#08#, 16#04#, 16#02#, 16#01#, -- x90
16#00#, 16#00#, 16#00#, 16#00#, 16#03#, 16#0c#, 16#30#, 16#c0#, 16#03#, 16#0c#, 16#30#, 16#c0#, 16#00#, 16#00#, 16#00#, 16#00#,
16#03#, 16#0c#, 16#30#, 16#c0#, 16#c0#, 16#30#, 16#0c#, 16#03#, 16#00#, 16#00#, 16#00#, 16#00#, 16#c0#, 16#30#, 16#0c#, 16#03#,
16#c0#, 16#30#, 16#0c#, 16#03#, 16#00#, 16#00#, 16#00#, 16#00#, 16#c0#, 16#30#, 16#0c#, 16#03#, 16#03#, 16#0c#, 16#30#, 16#c0#,
16#10#, 16#10#, 16#20#, 16#20#, 16#40#, 16#40#, 16#80#, 16#80#, 16#01#, 16#01#, 16#02#, 16#02#, 16#04#, 16#04#, 16#08#, 16#08#, -- x98
16#81#, 16#81#, 16#42#, 16#42#, 16#24#, 16#24#, 16#18#, 16#18#, 16#80#, 16#80#, 16#40#, 16#40#, 16#20#, 16#20#, 16#10#, 16#10#,
16#08#, 16#08#, 16#04#, 16#04#, 16#02#, 16#02#, 16#01#, 16#01#, 16#18#, 16#18#, 16#24#, 16#24#, 16#42#, 16#42#, 16#81#, 16#81#,
16#ff#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#80#, 16#80#, 16#80#, 16#80#, 16#80#, 16#80#, 16#80#, 16#80#,
16#00#, 16#00#, 16#00#, 16#ff#, 16#ff#, 16#00#, 16#00#, 16#00#, 16#18#, 16#18#, 16#18#, 16#18#, 16#18#, 16#18#, 16#18#, 16#18#, -- xA0
16#18#, 16#18#, 16#18#, 16#ff#, 16#ff#, 16#00#, 16#00#, 16#00#, 16#18#, 16#18#, 16#18#, 16#1f#, 16#1f#, 16#18#, 16#18#, 16#18#,
16#00#, 16#00#, 16#00#, 16#ff#, 16#ff#, 16#18#, 16#18#, 16#18#, 16#18#, 16#18#, 16#18#, 16#f8#, 16#f8#, 16#18#, 16#18#, 16#18#,
16#18#, 16#18#, 16#18#, 16#ff#, 16#ff#, 16#18#, 16#18#, 16#18#, 16#18#, 16#18#, 16#18#, 16#1f#, 16#1f#, 16#00#, 16#00#, 16#00#,
16#00#, 16#00#, 16#00#, 16#1f#, 16#1f#, 16#18#, 16#18#, 16#18#, 16#00#, 16#00#, 16#00#, 16#f8#, 16#f8#, 16#18#, 16#18#, 16#18#, -- xA8
16#18#, 16#18#, 16#18#, 16#f8#, 16#f8#, 16#00#, 16#00#, 16#00#, 16#80#, 16#80#, 16#80#, 16#40#, 16#40#, 16#20#, 16#18#, 16#07#,
16#01#, 16#01#, 16#01#, 16#02#, 16#02#, 16#04#, 16#18#, 16#e0#, 16#e0#, 16#18#, 16#04#, 16#02#, 16#02#, 16#01#, 16#01#, 16#01#,
16#07#, 16#18#, 16#20#, 16#40#, 16#40#, 16#80#, 16#80#, 16#80#, 16#81#, 16#42#, 16#24#, 16#18#, 16#18#, 16#24#, 16#42#, 16#81#,
16#f0#, 16#f0#, 16#f0#, 16#f0#, 16#00#, 16#00#, 16#00#, 16#00#, 16#0f#, 16#0f#, 16#0f#, 16#0f#, 16#00#, 16#00#, 16#00#, 16#00#, -- xB0
16#00#, 16#00#, 16#00#, 16#00#, 16#0f#, 16#0f#, 16#0f#, 16#0f#, 16#00#, 16#00#, 16#00#, 16#00#, 16#f0#, 16#f0#, 16#f0#, 16#f0#,
16#f0#, 16#f0#, 16#f0#, 16#f0#, 16#f0#, 16#f0#, 16#f0#, 16#f0#, 16#0f#, 16#0f#, 16#0f#, 16#0f#, 16#0f#, 16#0f#, 16#0f#, 16#0f#,
16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#ff#, 16#ff#, 16#ff#, 16#ff#,
16#f0#, 16#f0#, 16#f0#, 16#f0#, 16#0f#, 16#0f#, 16#0f#, 16#0f#, 16#0f#, 16#0f#, 16#0f#, 16#0f#, 16#f0#, 16#f0#, 16#f0#, 16#f0#, -- xB8
16#0f#, 16#0f#, 16#0f#, 16#0f#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#f0#, 16#f0#, 16#f0#, 16#f0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#,
16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#f0#, 16#f0#, 16#f0#, 16#f0#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#0f#, 16#0f#, 16#0f#, 16#0f#,
16#01#, 16#03#, 16#07#, 16#0f#, 16#1f#, 16#3f#, 16#7f#, 16#ff#, 16#ff#, 16#7f#, 16#3f#, 16#1f#, 16#0f#, 16#07#, 16#03#, 16#01#,
16#01#, 16#01#, 16#01#, 16#01#, 16#01#, 16#01#, 16#01#, 16#01#, 16#ff#, 16#80#, 16#80#, 16#80#, 16#80#, 16#80#, 16#80#, 16#80#, -- xC0
16#ff#, 16#80#, 16#80#, 16#9c#, 16#9c#, 16#9c#, 16#80#, 16#80#, 16#ff#, 16#ff#, 16#ff#, 16#e3#, 16#e3#, 16#e3#, 16#ff#, 16#ff#,
16#18#, 16#3c#, 16#7e#, 16#3c#, 16#18#, 16#3c#, 16#7e#, 16#ff#, 16#ff#, 16#00#, 16#ff#, 16#00#, 16#ff#, 16#00#, 16#ff#, 16#00#,
16#aa#, 16#aa#, 16#aa#, 16#aa#, 16#aa#, 16#aa#, 16#aa#, 16#aa#, 16#55#, 16#aa#, 16#55#, 16#aa#, 16#55#, 16#aa#, 16#55#, 16#aa#,
16#01#, 16#01#, 16#01#, 16#01#, 16#01#, 16#01#, 16#01#, 16#ff#, 16#00#, 16#10#, 16#38#, 16#7c#, 16#fe#, 16#7c#, 16#38#, 16#10#, -- xC8
16#38#, 16#10#, 16#92#, 16#fe#, 16#92#, 16#10#, 16#38#, 16#7c#, 16#00#, 16#6c#, 16#fe#, 16#fe#, 16#fe#, 16#7c#, 16#38#, 16#10#,
16#10#, 16#38#, 16#7c#, 16#fe#, 16#fe#, 16#7c#, 16#10#, 16#7c#, 16#e7#, 16#e7#, 16#42#, 16#ff#, 16#ff#, 16#42#, 16#e7#, 16#e7#,
16#db#, 16#ff#, 16#db#, 16#18#, 16#18#, 16#db#, 16#ff#, 16#db#, 16#3c#, 16#7e#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#7e#, 16#3c#,
16#c0#, 16#c0#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#30#, 16#30#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, -- xD0
16#0c#, 16#0c#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#03#, 16#03#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#,
16#00#, 16#00#, 16#c0#, 16#c0#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#30#, 16#30#, 16#00#, 16#00#, 16#00#, 16#00#,
16#00#, 16#00#, 16#0c#, 16#0c#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#03#, 16#03#, 16#00#, 16#00#, 16#00#, 16#00#,
16#00#, 16#00#, 16#00#, 16#00#, 16#c0#, 16#c0#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#30#, 16#30#, 16#00#, 16#00#, -- xD8
16#00#, 16#00#, 16#00#, 16#00#, 16#0c#, 16#0c#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#03#, 16#03#, 16#00#, 16#00#,
16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#c0#, 16#c0#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#30#, 16#30#,
16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#0c#, 16#0c#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#03#, 16#03#,
16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#0f#, 16#0f#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#3f#, 16#3f#, -- xE0
16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#ff#, 16#ff#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#fc#, 16#fc#,
16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#f0#, 16#f0#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#c0#, 16#c0#,
16#00#, 16#00#, 16#00#, 16#00#, 16#c0#, 16#c0#, 16#c0#, 16#c0#, 16#00#, 16#00#, 16#c0#, 16#c0#, 16#c0#, 16#c0#, 16#c0#, 16#c0#,
16#c0#, 16#c0#, 16#c0#, 16#c0#, 16#c0#, 16#c0#, 16#c0#, 16#c0#, 16#c0#, 16#c0#, 16#c0#, 16#c0#, 16#c0#, 16#c0#, 16#00#, 16#00#, -- xE8
16#c0#, 16#c0#, 16#c0#, 16#c0#, 16#00#, 16#00#, 16#00#, 16#00#, 16#c0#, 16#c0#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#,
16#f0#, 16#f0#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#fc#, 16#fc#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#,
16#ff#, 16#ff#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#3f#, 16#3f#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#,
16#0f#, 16#0f#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#03#, 16#03#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, -- xF0
16#03#, 16#03#, 16#03#, 16#03#, 16#00#, 16#00#, 16#00#, 16#00#, 16#03#, 16#03#, 16#03#, 16#03#, 16#03#, 16#03#, 16#00#, 16#00#,
16#03#, 16#03#, 16#03#, 16#03#, 16#03#, 16#03#, 16#03#, 16#03#, 16#00#, 16#00#, 16#03#, 16#03#, 16#03#, 16#03#, 16#03#, 16#03#,
16#00#, 16#00#, 16#00#, 16#00#, 16#03#, 16#03#, 16#03#, 16#03#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#03#, 16#03#,
16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#ff#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#ff#, 16#ff#, -- xF8
16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#ff#, 16#ff#, 16#ff#, 16#00#, 16#00#, 16#00#, 16#00#, 16#ff#, 16#ff#, 16#ff#, 16#ff#,
16#00#, 16#00#, 16#00#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#00#, 16#00#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#,
16#00#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#);
end package bm100_pkg;

