
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.bm100_pkg.all;                 -- character ROM type


entity charrom2 is
    port
    (
        clk         : in  std_logic;
        --
        addr_char_i : in  std_logic_vector(7 downto 0);
        addr_line_i : in  std_logic_vector(2 downto 0);
        --
        data_o      : out std_logic_vector(7 downto 0)
    );
end entity charrom2;


architecture rtl of charrom2 is

    constant rom_init_file : string := "../ROMs/ibm_zg+din.bin";

    -- function work with ModelSim (and Xilinx ISE) but not with Quartus 13.1!
    impure function init_crom( filename : string) return T_BM100_MEM is
        type charfile is file of character;
        file data_file  : charfile;
        variable rom    : T_BM100_MEM;
        variable c      : character;
    begin
        if filename'length = 0 then
            report init_crom'instance_name & " no filename given, ROM empty" severity warning;
            return rom;
        end if;

        file_open( data_file, filename, read_mode);
        for index in rom'range loop
            read( data_file, c);
            rom( index) := character'pos( c);
        end loop;
        file_close( data_file);

        return rom;
    end function init_crom;

    --signal crom_array : T_BM100_MEM := init_crom( rom_init_file);

    -- workaround for Quartus
    constant charrom2_init : T_BM100_MEM := (
        16#00#, 16#44#, 16#aa#, 16#aa#, 16#aa#, 16#aa#, 16#44#, 16#00#, -- 0
        16#40#, 16#a0#, 16#0c#, 16#12#, 16#1e#, 16#12#, 16#12#, 16#00#, -- 1
        16#40#, 16#a0#, 16#1c#, 16#12#, 16#1c#, 16#12#, 16#1c#, 16#00#, -- 2
        16#40#, 16#a0#, 16#0c#, 16#12#, 16#10#, 16#12#, 16#0c#, 16#00#, -- 3
        16#40#, 16#a0#, 16#1c#, 16#12#, 16#12#, 16#12#, 16#1c#, 16#00#, -- 4
        16#40#, 16#a0#, 16#1e#, 16#10#, 16#1c#, 16#10#, 16#1e#, 16#00#, -- 5
        16#40#, 16#a0#, 16#1e#, 16#10#, 16#1c#, 16#10#, 16#10#, 16#00#, -- 6
        16#40#, 16#a0#, 16#0c#, 16#12#, 16#10#, 16#16#, 16#0e#, 16#00#, -- 7
        16#40#, 16#a0#, 16#12#, 16#12#, 16#1e#, 16#12#, 16#12#, 16#00#, -- 8
        16#40#, 16#a0#, 16#0e#, 16#04#, 16#04#, 16#04#, 16#0e#, 16#00#, -- 9
        16#00#, 16#00#, 16#8e#, 16#88#, 16#8c#, 16#88#, 16#e8#, 16#00#, -- 10
        16#40#, 16#a0#, 16#12#, 16#14#, 16#18#, 16#14#, 16#12#, 16#00#, -- 11
        16#40#, 16#a0#, 16#10#, 16#10#, 16#10#, 16#10#, 16#1e#, 16#00#, -- 12
        16#00#, 16#00#, 16#6c#, 16#8a#, 16#8c#, 16#8a#, 16#6a#, 16#00#, -- 13
        16#40#, 16#a0#, 16#12#, 16#1a#, 16#16#, 16#12#, 16#12#, 16#00#, -- 14
        16#40#, 16#a0#, 16#0c#, 16#12#, 16#12#, 16#12#, 16#0c#, 16#00#, -- 15
        16#40#, 16#a0#, 16#1c#, 16#12#, 16#1c#, 16#10#, 16#10#, 16#00#, -- 16
        16#40#, 16#a0#, 16#0c#, 16#12#, 16#12#, 16#14#, 16#0a#, 16#00#, -- 17
        16#40#, 16#a0#, 16#1c#, 16#12#, 16#1c#, 16#14#, 16#12#, 16#00#, -- 18
        16#40#, 16#a0#, 16#0e#, 16#10#, 16#0c#, 16#02#, 16#1c#, 16#00#, -- 19
        16#40#, 16#a0#, 16#0e#, 16#04#, 16#04#, 16#04#, 16#04#, 16#00#, -- 20
        16#40#, 16#a0#, 16#12#, 16#12#, 16#12#, 16#12#, 16#0c#, 16#00#, -- 21
        16#40#, 16#a0#, 16#11#, 16#11#, 16#11#, 16#0a#, 16#04#, 16#00#, -- 22
        16#40#, 16#a0#, 16#11#, 16#15#, 16#15#, 16#1b#, 16#11#, 16#00#, -- 23
        16#40#, 16#a0#, 16#11#, 16#0a#, 16#04#, 16#0a#, 16#11#, 16#00#, -- 24
        16#40#, 16#a0#, 16#11#, 16#11#, 16#0a#, 16#04#, 16#04#, 16#00#, -- 25
        16#40#, 16#a0#, 16#1e#, 16#02#, 16#04#, 16#08#, 16#1e#, 16#00#, -- 26
        16#00#, 16#00#, 16#db#, 16#92#, 16#ca#, 16#8a#, 16#db#, 16#00#, -- 27
        16#48#, 16#a8#, 16#08#, 16#08#, 16#08#, 16#08#, 16#08#, 16#00#, -- 28
        16#40#, 16#a0#, 16#0c#, 16#04#, 16#06#, 16#04#, 16#0c#, 16#00#, -- 29
        16#00#, 16#00#, 16#94#, 16#d4#, 16#b4#, 16#94#, 16#96#, 16#00#, -- 30
        16#00#, 16#00#, 16#2e#, 16#68#, 16#2c#, 16#28#, 16#28#, 16#00#, -- 31
        16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, -- 32
        16#10#, 16#10#, 16#10#, 16#10#, 16#00#, 16#00#, 16#10#, 16#00#, -- 33
        16#28#, 16#28#, 16#28#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, -- 34
        16#24#, 16#7e#, 16#24#, 16#24#, 16#24#, 16#7e#, 16#24#, 16#00#, -- 35
        16#10#, 16#3c#, 16#50#, 16#38#, 16#14#, 16#78#, 16#10#, 16#00#, -- 36
        16#60#, 16#64#, 16#08#, 16#10#, 16#20#, 16#4c#, 16#0c#, 16#00#, -- 37
        16#10#, 16#28#, 16#28#, 16#30#, 16#54#, 16#48#, 16#34#, 16#00#, -- 38
        16#10#, 16#10#, 16#20#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, -- 39
        16#08#, 16#10#, 16#20#, 16#20#, 16#20#, 16#10#, 16#08#, 16#00#, -- 40
        16#20#, 16#10#, 16#08#, 16#08#, 16#08#, 16#10#, 16#20#, 16#00#, -- 41
        16#00#, 16#10#, 16#54#, 16#38#, 16#54#, 16#10#, 16#00#, 16#00#, -- 42
        16#00#, 16#10#, 16#10#, 16#7c#, 16#10#, 16#10#, 16#00#, 16#00#, -- 43
        16#00#, 16#00#, 16#00#, 16#00#, 16#10#, 16#10#, 16#20#, 16#00#, -- 44
        16#00#, 16#00#, 16#00#, 16#7c#, 16#00#, 16#00#, 16#00#, 16#00#, -- 45
        16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#30#, 16#30#, 16#00#, -- 46
        16#00#, 16#04#, 16#08#, 16#10#, 16#20#, 16#40#, 16#00#, 16#00#, -- 47
        16#38#, 16#44#, 16#4c#, 16#54#, 16#64#, 16#44#, 16#38#, 16#00#, -- 48
        16#10#, 16#30#, 16#10#, 16#10#, 16#10#, 16#10#, 16#38#, 16#00#, -- 49
        16#38#, 16#44#, 16#04#, 16#08#, 16#10#, 16#20#, 16#7c#, 16#00#, -- 50
        16#7c#, 16#08#, 16#10#, 16#08#, 16#04#, 16#44#, 16#38#, 16#00#, -- 51
        16#08#, 16#18#, 16#28#, 16#48#, 16#7c#, 16#08#, 16#08#, 16#00#, -- 52
        16#7c#, 16#40#, 16#78#, 16#04#, 16#04#, 16#44#, 16#38#, 16#00#, -- 53
        16#18#, 16#20#, 16#40#, 16#78#, 16#44#, 16#44#, 16#38#, 16#00#, -- 54
        16#7c#, 16#04#, 16#08#, 16#10#, 16#20#, 16#20#, 16#20#, 16#00#, -- 55
        16#38#, 16#44#, 16#44#, 16#38#, 16#44#, 16#44#, 16#38#, 16#00#, -- 56
        16#38#, 16#44#, 16#44#, 16#3c#, 16#04#, 16#08#, 16#30#, 16#00#, -- 57
        16#00#, 16#30#, 16#30#, 16#00#, 16#30#, 16#30#, 16#00#, 16#00#, -- 58
        16#00#, 16#00#, 16#10#, 16#00#, 16#10#, 16#10#, 16#20#, 16#00#, -- 59
        16#08#, 16#10#, 16#20#, 16#40#, 16#20#, 16#10#, 16#08#, 16#00#, -- 60
        16#00#, 16#00#, 16#7c#, 16#00#, 16#7c#, 16#00#, 16#00#, 16#00#, -- 61
        16#20#, 16#10#, 16#08#, 16#04#, 16#08#, 16#10#, 16#20#, 16#00#, -- 62
        16#38#, 16#44#, 16#04#, 16#08#, 16#10#, 16#00#, 16#10#, 16#00#, -- 63
        16#38#, 16#44#, 16#5c#, 16#54#, 16#5c#, 16#40#, 16#3c#, 16#00#, -- 64
        16#38#, 16#44#, 16#44#, 16#7c#, 16#44#, 16#44#, 16#44#, 16#00#, -- 65
        16#78#, 16#24#, 16#24#, 16#38#, 16#24#, 16#24#, 16#78#, 16#00#, -- 66
        16#38#, 16#44#, 16#40#, 16#40#, 16#40#, 16#44#, 16#38#, 16#00#, -- 67
        16#78#, 16#24#, 16#24#, 16#24#, 16#24#, 16#24#, 16#78#, 16#00#, -- 68
        16#7c#, 16#40#, 16#40#, 16#78#, 16#40#, 16#40#, 16#7c#, 16#00#, -- 69
        16#7c#, 16#40#, 16#40#, 16#78#, 16#40#, 16#40#, 16#40#, 16#00#, -- 70
        16#38#, 16#44#, 16#40#, 16#40#, 16#4c#, 16#44#, 16#3c#, 16#00#, -- 71
        16#44#, 16#44#, 16#44#, 16#7c#, 16#44#, 16#44#, 16#44#, 16#00#, -- 72
        16#38#, 16#10#, 16#10#, 16#10#, 16#10#, 16#10#, 16#38#, 16#00#, -- 73
        16#1c#, 16#08#, 16#08#, 16#08#, 16#08#, 16#48#, 16#30#, 16#00#, -- 74
        16#44#, 16#48#, 16#50#, 16#60#, 16#50#, 16#48#, 16#44#, 16#00#, -- 75
        16#40#, 16#40#, 16#40#, 16#40#, 16#40#, 16#40#, 16#7c#, 16#00#, -- 76
        16#44#, 16#6c#, 16#54#, 16#54#, 16#44#, 16#44#, 16#44#, 16#00#, -- 77
        16#44#, 16#44#, 16#64#, 16#54#, 16#4c#, 16#44#, 16#44#, 16#00#, -- 78
        16#38#, 16#44#, 16#44#, 16#44#, 16#44#, 16#44#, 16#38#, 16#00#, -- 79
        16#78#, 16#44#, 16#44#, 16#78#, 16#40#, 16#40#, 16#40#, 16#00#, -- 80
        16#38#, 16#44#, 16#44#, 16#44#, 16#54#, 16#48#, 16#34#, 16#00#, -- 81
        16#78#, 16#44#, 16#44#, 16#78#, 16#50#, 16#48#, 16#44#, 16#00#, -- 82
        16#3c#, 16#40#, 16#40#, 16#38#, 16#04#, 16#04#, 16#78#, 16#00#, -- 83
        16#7c#, 16#10#, 16#10#, 16#10#, 16#10#, 16#10#, 16#10#, 16#00#, -- 84
        16#44#, 16#44#, 16#44#, 16#44#, 16#44#, 16#44#, 16#38#, 16#00#, -- 85
        16#44#, 16#44#, 16#44#, 16#44#, 16#44#, 16#28#, 16#10#, 16#00#, -- 86
        16#44#, 16#44#, 16#44#, 16#54#, 16#54#, 16#6c#, 16#44#, 16#00#, -- 87
        16#44#, 16#44#, 16#28#, 16#10#, 16#28#, 16#44#, 16#44#, 16#00#, -- 88
        16#44#, 16#44#, 16#44#, 16#28#, 16#10#, 16#10#, 16#10#, 16#00#, -- 89
        16#7c#, 16#04#, 16#08#, 16#10#, 16#20#, 16#40#, 16#7c#, 16#00#, -- 90
        16#44#, 16#38#, 16#44#, 16#44#, 16#7c#, 16#44#, 16#44#, 16#00#, -- 91
        16#44#, 16#38#, 16#44#, 16#44#, 16#44#, 16#44#, 16#38#, 16#00#, -- 92
        16#44#, 16#00#, 16#44#, 16#44#, 16#44#, 16#44#, 16#38#, 16#00#, -- 93
        16#10#, 16#28#, 16#44#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, -- 94
        16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#7e#, 16#00#, -- 95
        16#00#, 16#20#, 16#10#, 16#08#, 16#00#, 16#00#, 16#00#, 16#00#, -- 96
        16#00#, 16#00#, 16#34#, 16#4c#, 16#44#, 16#44#, 16#3a#, 16#00#, -- 97
        16#40#, 16#40#, 16#58#, 16#64#, 16#44#, 16#44#, 16#78#, 16#00#, -- 98
        16#00#, 16#00#, 16#38#, 16#44#, 16#40#, 16#44#, 16#38#, 16#00#, -- 99
        16#04#, 16#04#, 16#34#, 16#4c#, 16#44#, 16#44#, 16#3a#, 16#00#, -- 100
        16#00#, 16#00#, 16#38#, 16#44#, 16#7c#, 16#40#, 16#38#, 16#00#, -- 101
        16#08#, 16#10#, 16#38#, 16#10#, 16#10#, 16#10#, 16#10#, 16#00#, -- 102
        16#00#, 16#00#, 16#34#, 16#4c#, 16#44#, 16#3c#, 16#04#, 16#38#, -- 103
        16#40#, 16#40#, 16#58#, 16#64#, 16#44#, 16#44#, 16#44#, 16#00#, -- 104
        16#10#, 16#00#, 16#10#, 16#10#, 16#10#, 16#10#, 16#08#, 16#00#, -- 105
        16#10#, 16#00#, 16#10#, 16#10#, 16#10#, 16#10#, 16#10#, 16#20#, -- 106
        16#40#, 16#40#, 16#48#, 16#50#, 16#70#, 16#48#, 16#44#, 16#00#, -- 107
        16#10#, 16#10#, 16#10#, 16#10#, 16#10#, 16#10#, 16#08#, 16#00#, -- 108
        16#00#, 16#00#, 16#68#, 16#54#, 16#54#, 16#54#, 16#54#, 16#00#, -- 109
        16#00#, 16#00#, 16#58#, 16#64#, 16#44#, 16#44#, 16#44#, 16#00#, -- 110
        16#00#, 16#00#, 16#38#, 16#44#, 16#44#, 16#44#, 16#38#, 16#00#, -- 111
        16#00#, 16#00#, 16#58#, 16#64#, 16#44#, 16#78#, 16#40#, 16#40#, -- 112
        16#00#, 16#00#, 16#34#, 16#4c#, 16#44#, 16#3c#, 16#04#, 16#04#, -- 113
        16#00#, 16#00#, 16#58#, 16#64#, 16#40#, 16#40#, 16#40#, 16#00#, -- 114
        16#00#, 16#00#, 16#38#, 16#40#, 16#38#, 16#04#, 16#78#, 16#00#, -- 115
        16#10#, 16#10#, 16#38#, 16#10#, 16#10#, 16#10#, 16#08#, 16#00#, -- 116
        16#00#, 16#00#, 16#44#, 16#44#, 16#44#, 16#4c#, 16#34#, 16#00#, -- 117
        16#00#, 16#00#, 16#44#, 16#44#, 16#44#, 16#28#, 16#10#, 16#00#, -- 118
        16#00#, 16#00#, 16#54#, 16#54#, 16#54#, 16#54#, 16#28#, 16#00#, -- 119
        16#00#, 16#00#, 16#44#, 16#28#, 16#10#, 16#28#, 16#44#, 16#00#, -- 120
        16#00#, 16#00#, 16#44#, 16#44#, 16#44#, 16#3c#, 16#04#, 16#38#, -- 121
        16#00#, 16#00#, 16#7c#, 16#08#, 16#10#, 16#20#, 16#7c#, 16#00#, -- 122
        16#28#, 16#00#, 16#34#, 16#4c#, 16#44#, 16#44#, 16#3a#, 16#00#, -- 123
        16#28#, 16#00#, 16#38#, 16#44#, 16#44#, 16#44#, 16#38#, 16#00#, -- 124
        16#28#, 16#00#, 16#44#, 16#44#, 16#44#, 16#4c#, 16#34#, 16#00#, -- 125
        16#18#, 16#24#, 16#24#, 16#28#, 16#24#, 16#34#, 16#28#, 16#00#, -- 126
        16#ff#, 16#cf#, 16#e7#, 16#f3#, 16#e7#, 16#cf#, 16#ff#, 16#00#, -- 127
        16#38#, 16#44#, 16#40#, 16#40#, 16#44#, 16#38#, 16#08#, 16#30#, -- 128
        16#28#, 16#00#, 16#44#, 16#44#, 16#44#, 16#44#, 16#3a#, 16#00#, -- 129
        16#08#, 16#10#, 16#38#, 16#44#, 16#7c#, 16#40#, 16#38#, 16#00#, -- 130
        16#38#, 16#44#, 16#38#, 16#04#, 16#3c#, 16#44#, 16#3a#, 16#00#, -- 131
        16#28#, 16#00#, 16#38#, 16#04#, 16#3c#, 16#44#, 16#3a#, 16#00#, -- 132
        16#20#, 16#10#, 16#38#, 16#04#, 16#3c#, 16#44#, 16#3a#, 16#00#, -- 133
        16#10#, 16#00#, 16#38#, 16#04#, 16#3c#, 16#44#, 16#3a#, 16#00#, -- 134
        16#00#, 16#00#, 16#38#, 16#44#, 16#40#, 16#44#, 16#38#, 16#08#, -- 135
        16#38#, 16#44#, 16#38#, 16#44#, 16#7c#, 16#40#, 16#38#, 16#00#, -- 136
        16#28#, 16#00#, 16#38#, 16#44#, 16#7c#, 16#40#, 16#38#, 16#00#, -- 137
        16#10#, 16#08#, 16#38#, 16#44#, 16#7c#, 16#40#, 16#38#, 16#00#, -- 138
        16#28#, 16#00#, 16#10#, 16#10#, 16#10#, 16#10#, 16#08#, 16#00#, -- 139
        16#38#, 16#44#, 16#10#, 16#10#, 16#10#, 16#10#, 16#08#, 16#00#, -- 140
        16#10#, 16#08#, 16#10#, 16#10#, 16#10#, 16#10#, 16#08#, 16#00#, -- 141
        16#44#, 16#10#, 16#28#, 16#44#, 16#44#, 16#7c#, 16#44#, 16#00#, -- 142
        16#28#, 16#44#, 16#38#, 16#44#, 16#44#, 16#7c#, 16#44#, 16#00#, -- 143
        16#08#, 16#10#, 16#7c#, 16#40#, 16#78#, 16#40#, 16#7c#, 16#00#, -- 144
        16#00#, 16#00#, 16#6c#, 16#14#, 16#7c#, 16#50#, 16#6c#, 16#00#, -- 145
        16#1c#, 16#30#, 16#50#, 16#7c#, 16#50#, 16#50#, 16#5c#, 16#00#, -- 146
        16#38#, 16#44#, 16#00#, 16#38#, 16#44#, 16#44#, 16#38#, 16#00#, -- 147
        16#28#, 16#00#, 16#38#, 16#44#, 16#44#, 16#44#, 16#38#, 16#00#, -- 148
        16#10#, 16#08#, 16#38#, 16#44#, 16#44#, 16#44#, 16#38#, 16#00#, -- 149
        16#38#, 16#44#, 16#00#, 16#44#, 16#44#, 16#44#, 16#3a#, 16#00#, -- 150
        16#20#, 16#10#, 16#44#, 16#44#, 16#44#, 16#44#, 16#3a#, 16#00#, -- 151
        16#28#, 16#00#, 16#44#, 16#44#, 16#44#, 16#3c#, 16#04#, 16#38#, -- 152
        16#44#, 16#38#, 16#44#, 16#44#, 16#44#, 16#44#, 16#38#, 16#00#, -- 153
        16#44#, 16#00#, 16#44#, 16#44#, 16#44#, 16#44#, 16#38#, 16#00#, -- 154
        16#00#, 16#10#, 16#3c#, 16#50#, 16#50#, 16#3c#, 16#10#, 16#00#, -- 155
        16#18#, 16#24#, 16#20#, 16#70#, 16#20#, 16#20#, 16#7c#, 16#00#, -- 156
        16#44#, 16#28#, 16#7c#, 16#10#, 16#7c#, 16#10#, 16#10#, 16#00#, -- 157
        16#20#, 16#50#, 16#40#, 16#64#, 16#4e#, 16#44#, 16#46#, 16#00#, -- 158
        16#18#, 16#24#, 16#20#, 16#78#, 16#20#, 16#20#, 16#60#, 16#00#, -- 159
        16#10#, 16#20#, 16#38#, 16#04#, 16#3c#, 16#44#, 16#3a#, 16#00#, -- 160
        16#08#, 16#10#, 16#00#, 16#10#, 16#10#, 16#10#, 16#08#, 16#00#, -- 161
        16#08#, 16#10#, 16#38#, 16#44#, 16#44#, 16#44#, 16#38#, 16#00#, -- 162
        16#08#, 16#10#, 16#44#, 16#44#, 16#44#, 16#44#, 16#3a#, 16#00#, -- 163
        16#20#, 16#54#, 16#08#, 16#58#, 16#64#, 16#44#, 16#44#, 16#00#, -- 164
        16#20#, 16#54#, 16#08#, 16#64#, 16#54#, 16#4c#, 16#44#, 16#00#, -- 165
        16#38#, 16#04#, 16#3c#, 16#44#, 16#3a#, 16#00#, 16#7c#, 16#00#, -- 166
        16#58#, 16#44#, 16#44#, 16#44#, 16#58#, 16#00#, 16#7c#, 16#00#, -- 167
        16#10#, 16#00#, 16#10#, 16#20#, 16#44#, 16#44#, 16#38#, 16#00#, -- 168
        16#00#, 16#00#, 16#00#, 16#00#, 16#7e#, 16#40#, 16#40#, 16#00#, -- 169
        16#00#, 16#00#, 16#00#, 16#00#, 16#7e#, 16#02#, 16#02#, 16#00#, -- 170
        16#44#, 16#48#, 16#50#, 16#2c#, 16#52#, 16#04#, 16#0e#, 16#00#, -- 171
        16#44#, 16#48#, 16#50#, 16#2c#, 16#54#, 16#1e#, 16#04#, 16#00#, -- 172
        16#10#, 16#00#, 16#10#, 16#10#, 16#10#, 16#10#, 16#10#, 16#00#, -- 173
        16#00#, 16#00#, 16#12#, 16#24#, 16#48#, 16#24#, 16#12#, 16#00#, -- 174
        16#00#, 16#00#, 16#48#, 16#24#, 16#12#, 16#24#, 16#48#, 16#00#, -- 175
        16#55#, 16#00#, 16#55#, 16#00#, 16#55#, 16#00#, 16#55#, 16#00#, -- 176
        16#55#, 16#aa#, 16#55#, 16#aa#, 16#55#, 16#aa#, 16#55#, 16#aa#, -- 177
        16#aa#, 16#55#, 16#aa#, 16#55#, 16#aa#, 16#55#, 16#aa#, 16#55#, -- 178
        16#10#, 16#10#, 16#10#, 16#10#, 16#10#, 16#10#, 16#10#, 16#10#, -- 179
        16#10#, 16#10#, 16#10#, 16#10#, 16#f0#, 16#10#, 16#10#, 16#10#, -- 180
        16#10#, 16#10#, 16#f0#, 16#10#, 16#f0#, 16#10#, 16#10#, 16#10#, -- 181
        16#14#, 16#14#, 16#14#, 16#14#, 16#f4#, 16#14#, 16#14#, 16#14#, -- 182
        16#00#, 16#00#, 16#00#, 16#00#, 16#fc#, 16#14#, 16#14#, 16#14#, -- 183
        16#00#, 16#00#, 16#f0#, 16#10#, 16#f0#, 16#10#, 16#10#, 16#10#, -- 184
        16#14#, 16#14#, 16#f4#, 16#04#, 16#f4#, 16#14#, 16#14#, 16#14#, -- 185
        16#14#, 16#14#, 16#14#, 16#14#, 16#14#, 16#14#, 16#14#, 16#14#, -- 186
        16#00#, 16#00#, 16#fc#, 16#04#, 16#f4#, 16#14#, 16#14#, 16#14#, -- 187
        16#14#, 16#14#, 16#f4#, 16#04#, 16#fc#, 16#00#, 16#00#, 16#00#, -- 188
        16#14#, 16#14#, 16#14#, 16#14#, 16#fc#, 16#00#, 16#00#, 16#00#, -- 189
        16#10#, 16#10#, 16#f0#, 16#10#, 16#f0#, 16#00#, 16#00#, 16#00#, -- 190
        16#00#, 16#00#, 16#00#, 16#00#, 16#f0#, 16#10#, 16#10#, 16#10#, -- 191
        16#10#, 16#10#, 16#10#, 16#10#, 16#1f#, 16#00#, 16#00#, 16#00#, -- 192
        16#10#, 16#10#, 16#10#, 16#10#, 16#ff#, 16#00#, 16#00#, 16#00#, -- 193
        16#00#, 16#00#, 16#00#, 16#00#, 16#ff#, 16#10#, 16#10#, 16#10#, -- 194
        16#10#, 16#10#, 16#10#, 16#10#, 16#1f#, 16#10#, 16#10#, 16#10#, -- 195
        16#00#, 16#00#, 16#00#, 16#00#, 16#ff#, 16#00#, 16#00#, 16#00#, -- 196
        16#10#, 16#10#, 16#10#, 16#10#, 16#ff#, 16#10#, 16#10#, 16#10#, -- 197
        16#10#, 16#10#, 16#1f#, 16#10#, 16#1f#, 16#10#, 16#10#, 16#10#, -- 198
        16#14#, 16#14#, 16#14#, 16#14#, 16#17#, 16#14#, 16#14#, 16#14#, -- 199
        16#14#, 16#14#, 16#17#, 16#10#, 16#1f#, 16#00#, 16#00#, 16#00#, -- 200
        16#00#, 16#00#, 16#1f#, 16#10#, 16#17#, 16#14#, 16#14#, 16#14#, -- 201
        16#14#, 16#14#, 16#f7#, 16#00#, 16#ff#, 16#00#, 16#00#, 16#00#, -- 202
        16#00#, 16#00#, 16#ff#, 16#00#, 16#f7#, 16#14#, 16#14#, 16#14#, -- 203
        16#14#, 16#14#, 16#17#, 16#10#, 16#17#, 16#14#, 16#14#, 16#14#, -- 204
        16#00#, 16#00#, 16#ff#, 16#00#, 16#ff#, 16#00#, 16#00#, 16#00#, -- 205
        16#14#, 16#14#, 16#f7#, 16#00#, 16#f7#, 16#14#, 16#14#, 16#14#, -- 206
        16#10#, 16#10#, 16#ff#, 16#00#, 16#ff#, 16#00#, 16#00#, 16#00#, -- 207
        16#14#, 16#14#, 16#14#, 16#14#, 16#ff#, 16#00#, 16#00#, 16#00#, -- 208
        16#00#, 16#00#, 16#ff#, 16#00#, 16#ff#, 16#10#, 16#10#, 16#10#, -- 209
        16#00#, 16#00#, 16#00#, 16#00#, 16#ff#, 16#14#, 16#14#, 16#14#, -- 210
        16#14#, 16#14#, 16#14#, 16#14#, 16#1f#, 16#00#, 16#00#, 16#00#, -- 211
        16#10#, 16#10#, 16#1f#, 16#10#, 16#1f#, 16#00#, 16#00#, 16#00#, -- 212
        16#00#, 16#00#, 16#1f#, 16#10#, 16#1f#, 16#10#, 16#10#, 16#10#, -- 213
        16#00#, 16#00#, 16#00#, 16#00#, 16#1f#, 16#14#, 16#14#, 16#14#, -- 214
        16#14#, 16#14#, 16#14#, 16#14#, 16#f7#, 16#14#, 16#14#, 16#14#, -- 215
        16#10#, 16#10#, 16#ff#, 16#00#, 16#ff#, 16#10#, 16#10#, 16#10#, -- 216
        16#10#, 16#10#, 16#10#, 16#10#, 16#f0#, 16#00#, 16#00#, 16#00#, -- 217
        16#00#, 16#00#, 16#00#, 16#00#, 16#1f#, 16#10#, 16#10#, 16#10#, -- 218
        16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, -- 219
        16#00#, 16#00#, 16#00#, 16#00#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, -- 220
        16#f0#, 16#f0#, 16#f0#, 16#f0#, 16#f0#, 16#f0#, 16#f0#, 16#f0#, -- 221
        16#0f#, 16#0f#, 16#0f#, 16#0f#, 16#0f#, 16#0f#, 16#0f#, 16#0f#, -- 222
        16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#00#, 16#00#, 16#00#, 16#00#, -- 223
        16#00#, 16#00#, 16#02#, 16#74#, 16#48#, 16#58#, 16#66#, 16#00#, -- 224
        16#18#, 16#24#, 16#24#, 16#28#, 16#24#, 16#34#, 16#28#, 16#00#, -- 225
        16#7c#, 16#44#, 16#40#, 16#40#, 16#40#, 16#40#, 16#40#, 16#00#, -- 226
        16#00#, 16#00#, 16#7c#, 16#28#, 16#28#, 16#28#, 16#4c#, 16#00#, -- 227
        16#7e#, 16#22#, 16#10#, 16#08#, 16#10#, 16#22#, 16#7e#, 16#00#, -- 228
        16#00#, 16#02#, 16#3c#, 16#48#, 16#48#, 16#48#, 16#30#, 16#00#, -- 229
        16#00#, 16#00#, 16#24#, 16#24#, 16#24#, 16#24#, 16#5c#, 16#80#, -- 230
        16#00#, 16#00#, 16#3e#, 16#80#, 16#10#, 16#10#, 16#18#, 16#00#, -- 231
        16#38#, 16#10#, 16#38#, 16#54#, 16#38#, 16#10#, 16#38#, 16#00#, -- 232
        16#38#, 16#44#, 16#44#, 16#7c#, 16#44#, 16#44#, 16#38#, 16#00#, -- 233
        16#38#, 16#44#, 16#44#, 16#44#, 16#28#, 16#28#, 16#6c#, 16#00#, -- 234
        16#04#, 16#08#, 16#08#, 16#38#, 16#44#, 16#44#, 16#38#, 16#00#, -- 235
        16#00#, 16#6c#, 16#92#, 16#92#, 16#92#, 16#6c#, 16#00#, 16#00#, -- 236
        16#02#, 16#3c#, 16#4c#, 16#54#, 16#64#, 16#78#, 16#80#, 16#00#, -- 237
        16#1e#, 16#20#, 16#40#, 16#7e#, 16#40#, 16#20#, 16#1e#, 16#00#, -- 238
        16#38#, 16#44#, 16#44#, 16#44#, 16#44#, 16#44#, 16#44#, 16#00#, -- 239
        16#00#, 16#00#, 16#7e#, 16#00#, 16#7e#, 16#00#, 16#7e#, 16#00#, -- 240
        16#10#, 16#10#, 16#7c#, 16#10#, 16#10#, 16#00#, 16#7c#, 16#00#, -- 241
        16#20#, 16#10#, 16#08#, 16#10#, 16#20#, 16#00#, 16#7c#, 16#00#, -- 242
        16#08#, 16#10#, 16#20#, 16#10#, 16#08#, 16#00#, 16#7c#, 16#00#, -- 243
        16#08#, 16#14#, 16#10#, 16#10#, 16#10#, 16#10#, 16#10#, 16#10#, -- 244
        16#10#, 16#10#, 16#10#, 16#10#, 16#10#, 16#10#, 16#50#, 16#20#, -- 245
        16#30#, 16#30#, 16#00#, 16#fc#, 16#00#, 16#30#, 16#30#, 16#00#, -- 246
        16#00#, 16#20#, 16#54#, 16#08#, 16#20#, 16#54#, 16#08#, 16#00#, -- 247
        16#18#, 16#24#, 16#24#, 16#18#, 16#00#, 16#00#, 16#00#, 16#00#, -- 248
        16#00#, 16#18#, 16#3c#, 16#18#, 16#00#, 16#00#, 16#00#, 16#00#, -- 249
        16#00#, 16#18#, 16#18#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, -- 250
        16#07#, 16#04#, 16#04#, 16#64#, 16#14#, 16#0c#, 16#0c#, 16#04#, -- 251
        16#28#, 16#34#, 16#24#, 16#24#, 16#24#, 16#00#, 16#00#, 16#00#, -- 252
        16#18#, 16#24#, 16#08#, 16#10#, 16#3c#, 16#00#, 16#00#, 16#00#, -- 253
        16#00#, 16#00#, 16#38#, 16#38#, 16#38#, 16#38#, 16#00#, 16#00#, -- 254
        16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#81#, 16#ff#, 16#ff#  -- 255
    );

    signal crom_array : T_BM100_MEM := charrom2_init;
    signal crom_index : natural;


begin

    crom_index <= to_integer( unsigned( addr_char_i & addr_line_i));
  
    process
    begin
        wait until rising_edge( clk);
        data_o <= std_logic_vector( to_unsigned( crom_array( crom_index), 8));
    end process;

end architecture rtl;
