------------------------------------------------------------------------
-- vga_controller_800_600.vhd
------------------------------------------------------------------------
-- Author : Ulrich Zolt�n
--          Copyright 2006 Digilent, Inc.
--
-- following things where changed by Bert Lange 2018:
--   - if rising_edge --> wait until rising_edge
--   - binary init values to readable integers
--   - add xFACTOR function
--   - change horizontal vales to use 60 MHz pixel clock for 800x600 timing
--     the 1200 pixels where combined later to 600 or 400 pixels
------------------------------------------------------------------------
--
--  the original Z1013 has 32x32 char video mode
--  with peters addition 
--
--   modes  chars pixels   *x    x   2*y percent of width
--   -----  ----- ------- ---- ---- ---- ----------------
--   32x32  32x32 256x256  3    768  512  64
--   64x16  64x32 512x256  2   1024  512  85
--
------------------------------------------------------------------------
-- Software version : Xilinx ISE 7.1.04i
--                    WebPack
-- Device	        : 3s200ft256-4
------------------------------------------------------------------------
-- This file contains the logic to generate the synchronization signals,
-- horizontal and vertical pixel counter and video disable signal
-- for the 800x600@60Hz resolution.
------------------------------------------------------------------------
--  Behavioral description
------------------------------------------------------------------------
-- Please read the following article on the web regarding the
-- vga video timings:
-- http://www.epanorama.net/documents/pc/vga_timing.html

-- This module generates the video synch pulses for the monitor to
-- enter 800x600@60Hz resolution state. It also provides horizontal
-- and vertical counters for the currently displayed pixel and a blank
-- signal that is active when the pixel is not inside the visible screen
-- and the color outputs should be reset to 0.

-- timing diagram for the horizontal synch signal (HS)
-- 0                         840    968          1056 (pixels)
-- _________________________|------|_________________
-- timing diagram for the vertical synch signal (VS)
-- 0                                  601    605  628 (lines)
-- __________________________________|------|________

-- The blank signal is delayed one pixel clock period (25ns) from where
-- the pixel leaves the visible screen, according to the counters, to
-- account for the pixel pipeline delay. This delay happens because
-- it takes time from when the counters indicate current pixel should
-- be displayed to when the color data actually arrives at the monitor
-- pins (memory read delays, synchronization delays).
------------------------------------------------------------------------
--  Port definitions
------------------------------------------------------------------------
-- rst               - global reset signal
-- pixel_clk         - input pin, from dcm_40MHz
--                   - the clock signal generated by a DCM that has
--                   - a frequency of 40MHz.
-- HS                - output pin, to monitor
--                   - horizontal synch pulse
-- VS                - output pin, to monitor
--                   - vertical synch pulse
-- hcount            - output pin, 11 bits, to clients
--                   - horizontal count of the currently displayed
--                   - pixel (even if not in visible area)
-- vcount            - output pin, 11 bits, to clients
--                   - vertical count of the currently active video
--                   - line (even if not in visible area)
-- blank             - output pin, to clients
--                   - active when pixel is not in visible area.
------------------------------------------------------------------------
-- Revision History:
-- 09/18/2006(UlrichZ): created
------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


-- the vga_controller_800_600 entity declaration
-- read above for behavioral description and port definitions.
entity vga_controller_800_600 is
port(
   rst         : in std_logic;
   pixel_clk   : in std_logic;
   --
   HS          : out std_logic;
   VS          : out std_logic;
   hcount      : out unsigned(10 downto 0);
   vcount      : out unsigned(10 downto 0);
   blank       : out std_logic
);
end entity vga_controller_800_600;


architecture Behavioral of vga_controller_800_600 is

------------------------------------------------------------------------
-- CONSTANTS
------------------------------------------------------------------------

-- factor for horizontal timing (pixel_clk/40MHz = 1.5)
function xFACTOR( x : integer) return integer is
begin
    return x + x / 2;
end function;

-- maximum value for the horizontal pixel counter
constant HMAX  : unsigned(10 downto 0) := to_unsigned( xFACTOR( 1056), 11); --"10000100000";

-- maximum value for the vertical pixel counter
constant VMAX  : unsigned(10 downto 0) := to_unsigned(  628, 11);           --"01001110100";

-- total number of visible columns
constant HLINES: unsigned(10 downto 0) := to_unsigned( xFACTOR( 800), 11);  --"01100100000";

-- value for the horizontal counter where front porch ends
constant HFP   : unsigned(10 downto 0) := to_unsigned( xFACTOR( 840), 11);  --"01101001000";

-- value for the horizontal counter where the synch pulse ends
constant HSP   : unsigned(10 downto 0) := to_unsigned( xFACTOR( 968), 11);  --"01111001000";

-- total number of visible lines
constant VLINES: unsigned(10 downto 0) := to_unsigned(  600, 11);           --"01001011000";

-- value for the vertical counter where the front porch ends
constant VFP   : unsigned(10 downto 0) := to_unsigned(  601, 11);           --"01001011001";

-- value for the vertical counter where the synch pulse ends
constant VSP   : unsigned(10 downto 0) := to_unsigned(  605, 11);           --"01001011101";

-- polarity of the horizontal and vertical synch pulse
-- only one polarity used, because for this resolution they coincide.
constant SPP   : std_logic := '1';

------------------------------------------------------------------------
-- SIGNALS
------------------------------------------------------------------------

-- horizontal and vertical counters
signal hcounter : unsigned(10 downto 0) := (others => '0');
signal vcounter : unsigned(10 downto 0) := (others => '0');

-- active when inside visible screen area.
signal video_enable: std_logic;

begin

   -- output horizontal and vertical counters
   hcount <= hcounter;
   vcount <= vcounter;

   -- blank is active when outside screen visible area
   -- color output should be blacked (put on 0) when blank in active
   -- blank is delayed one pixel clock period from the video_enable
   -- signal to account for the pixel pipeline delay.
   blank <= not video_enable when rising_edge(pixel_clk);

   -- increment horizontal counter at pixel_clk rate
   -- until HMAX is reached, then reset and keep counting
   h_count: process
   begin
      wait until rising_edge(pixel_clk);
      if(rst = '1') then
         hcounter <= (others => '0');
      elsif(hcounter = HMAX) then
         hcounter <= (others => '0');
      else
         hcounter <= hcounter + 1;
      end if;
   end process h_count;

   -- increment vertical counter when one line is finished
   -- (horizontal counter reached HMAX)
   -- until VMAX is reached, then reset and keep counting
   v_count: process
   begin
      wait until rising_edge(pixel_clk);
      if(rst = '1') then
         vcounter <= (others => '0');
      elsif(hcounter = HMAX) then
         if(vcounter = VMAX) then
            vcounter <= (others => '0');
         else
            vcounter <= vcounter + 1;
         end if;
      end if;
   end process v_count;

   -- generate horizontal synch pulse
   -- when horizontal counter is between where the
   -- front porch ends and the synch pulse ends.
   -- The HS is active (with polarity SPP) for a total of 128 pixels.
   do_hs: process
   begin
      wait until rising_edge(pixel_clk);
      if(hcounter >= HFP and hcounter < HSP) then
         HS <= not SPP;
      else
         HS <= SPP;
      end if;
   end process do_hs;

   -- generate vertical synch pulse
   -- when vertical counter is between where the
   -- front porch ends and the synch pulse ends.
   -- The VS is active (with polarity SPP) for a total of 4 video lines
   -- = 4*HMAX = 4224 pixels.
   do_vs: process
   begin
      wait until rising_edge(pixel_clk);
      if(vcounter >= VFP and vcounter < VSP) then
         VS <= not SPP;
      else
         VS <= SPP;
      end if;
   end process do_vs;
   
   -- enable video output when pixel is in visible area
   video_enable <= '1' when (hcounter < HLINES and vcounter < VLINES) else '0';

end Behavioral;
