----------------------------------------------------------------------------------
-- small 5x8 bitmap font (ASCII 32..127)
-- 
-- Copyright (c) 2017 by Bert Lange
-- https://github.com/boert/Z1013-mist
-- 
-- This source file is free software: you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published
-- by the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
-- 
-- This source file is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
-- 
-- You should have received a copy of the GNU General Public License
-- along with this program.  If not, see <http://www.gnu.org/licenses/>.
-- 
----------------------------------------------------------------------------------


package chars is

type chars_t is array(natural range <>) of integer;
constant chars_size       : natural := 10000;
constant chars : chars_t(0 to chars_size-1) := (
-- 
0,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- !
0,1,0,0,0,
0,1,0,0,0,
0,1,0,0,0,
0,1,0,0,0,
0,0,0,0,0,
0,1,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- "
0,0,0,0,0,
0,1,0,1,0,
0,1,0,1,0,
0,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- #
0,1,0,1,0,
0,1,0,1,0,
1,1,1,1,1,
0,1,0,1,0,
1,1,1,1,1,
0,1,0,1,0,
0,0,0,0,0,
0,0,0,0,0,
-- $
0,0,1,0,0,
0,1,1,1,0,
1,0,0,0,0,
0,1,1,1,0,
0,0,0,1,0,
0,1,1,1,0,
0,0,1,0,0,
0,0,0,0,0,
-- %
0,0,0,0,0,
0,1,0,1,0,
0,0,0,1,0,
0,0,1,0,0,
0,0,1,0,0,
0,1,0,0,0,
0,1,0,1,0,
0,0,0,0,0,
-- '
0,0,0,0,0,
0,1,0,0,0,
0,1,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- &
0,1,1,0,0,
1,0,0,0,0,
1,0,1,0,0,
0,1,0,0,0,
1,0,1,0,0,
0,1,0,1,0,
0,0,0,0,0,
0,0,0,0,0,
-- (
0,1,0,0,0,
1,0,0,0,0,
1,0,0,0,0,
1,0,0,0,0,
1,0,0,0,0,
0,1,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- )
1,0,0,0,0,
0,1,0,0,0,
0,1,0,0,0,
0,1,0,0,0,
0,1,0,0,0,
1,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- *
0,0,0,0,0,
1,0,0,1,0,
0,1,1,0,0,
1,1,1,1,0,
0,1,1,0,0,
1,0,0,1,0,
0,0,0,0,0,
0,0,0,0,0,
-- +
0,0,0,0,0,
0,0,1,0,0,
0,0,1,0,0,
1,1,1,1,1,
0,0,1,0,0,
0,0,1,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- ,
0,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
0,1,0,0,0,
1,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- -
0,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
1,1,1,1,1,
0,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- .
0,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
0,1,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- /
0,0,1,0,0,
0,0,1,0,0,
0,1,0,0,0,
0,1,0,0,0,
1,0,0,0,0,
1,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- 0
0,0,0,0,0,
0,1,1,0,0,
1,0,1,1,0,
1,0,0,1,0,
1,1,0,1,0,
0,1,1,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- 1
0,0,0,0,0,
0,0,1,1,0,
0,1,0,1,0,
0,0,0,1,0,
0,0,0,1,0,
0,0,0,1,0,
0,0,0,0,0,
0,0,0,0,0,
-- 2
0,0,0,0,0,
0,1,1,0,0,
1,0,0,1,0,
0,0,1,0,0,
0,1,0,0,0,
1,1,1,1,0,
0,0,0,0,0,
0,0,0,0,0,
-- 3
0,0,0,0,0,
0,1,1,0,0,
1,0,0,1,0,
0,0,1,0,0,
0,0,0,1,0,
1,0,0,1,0,
0,1,1,0,0,
0,0,0,0,0,
-- 4
0,0,0,0,0,
1,0,0,0,0,
1,0,0,0,0,
1,0,1,0,0,
1,1,1,1,0,
0,0,1,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- 5
0,0,0,0,0,
1,1,1,1,0,
1,0,0,0,0,
1,1,1,0,0,
0,0,0,1,0,
1,1,1,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- 6
0,0,0,0,0,
0,1,1,0,0,
1,0,0,1,0,
1,1,1,0,0,
1,0,0,1,0,
0,1,1,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- 7
0,0,0,0,0,
1,1,1,1,0,
0,0,0,1,0,
0,0,1,0,0,
0,0,1,0,0,
0,1,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- 8
0,0,0,0,0,
0,1,1,0,0,
1,0,0,1,0,
0,1,1,0,0,
1,0,0,1,0,
0,1,1,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- 9
0,0,0,0,0,
0,1,1,0,0,
1,0,0,1,0,
0,1,1,0,0,
0,0,0,1,0,
0,1,1,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- :
0,0,0,0,0,
0,0,0,0,0,
0,1,0,0,0,
0,0,0,0,0,
0,1,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- ;
0,0,0,0,0,
0,0,0,0,0,
0,1,0,0,0,
0,0,0,0,0,
0,1,0,0,0,
1,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- <
0,0,0,0,0,
0,0,1,0,0,
0,1,0,0,0,
1,0,0,0,0,
0,1,0,0,0,
0,0,1,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- =
0,0,0,0,0,
0,0,0,0,0,
1,1,1,1,0,
0,0,0,0,0,
1,1,1,1,0,
0,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- >
0,0,0,0,0,
0,1,0,0,0,
0,0,1,0,0,
0,0,0,1,0,
0,0,1,0,0,
0,1,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- ?
0,1,1,0,0,
1,0,0,1,0,
0,0,0,1,0,
0,0,1,0,0,
0,0,1,0,0,
0,0,0,0,0,
0,0,1,0,0,
0,0,0,0,0,
-- @
0,0,0,0,0,
0,1,1,0,0,
1,0,0,1,0,
1,0,1,1,0,
1,0,1,1,0,
0,1,1,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- A
0,1,1,0,0,
1,0,0,1,0,
1,0,0,1,0,
1,1,1,1,0,
1,0,0,1,0,
1,0,0,1,0,
0,0,0,0,0,
0,0,0,0,0,
-- B
1,1,1,0,0,
1,0,0,1,0,
1,1,1,0,0,
1,0,0,1,0,
1,0,0,1,0,
1,1,1,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- C
0,1,1,0,0,
1,0,0,1,0,
1,0,0,0,0,
1,0,0,0,0,
1,0,0,1,0,
0,1,1,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- D
1,1,1,0,0,
1,0,0,1,0,
1,0,0,1,0,
1,0,0,1,0,
1,0,0,1,0,
1,1,1,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- E
1,1,1,1,0,
1,0,0,0,0,
1,1,1,0,0,
1,0,0,0,0,
1,0,0,0,0,
1,1,1,1,0,
0,0,0,0,0,
0,0,0,0,0,
-- F
1,1,1,1,0,
1,0,0,0,0,
1,1,1,0,0,
1,0,0,0,0,
1,0,0,0,0,
1,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- G
0,1,1,0,0,
1,0,0,1,0,
1,0,0,0,0,
1,0,1,1,0,
1,0,0,1,0,
0,1,1,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- H
1,0,0,1,0,
1,0,0,1,0,
1,1,1,1,0,
1,0,0,1,0,
1,0,0,1,0,
1,0,0,1,0,
0,0,0,0,0,
0,0,0,0,0,
-- I
1,1,1,0,0,
0,1,0,0,0,
0,1,0,0,0,
0,1,0,0,0,
0,1,0,0,0,
1,1,1,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- J
0,1,1,1,0,
0,0,0,1,0,
0,0,0,1,0,
0,0,0,1,0,
1,0,0,1,0,
0,1,1,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- K
1,0,0,1,0,
1,0,1,0,0,
1,1,0,0,0,
1,1,0,0,0,
1,0,1,0,0,
1,0,0,1,0,
0,0,0,0,0,
0,0,0,0,0,
-- L
1,0,0,0,0,
1,0,0,0,0,
1,0,0,0,0,
1,0,0,0,0,
1,0,0,1,0,
1,1,1,1,0,
0,0,0,0,0,
0,0,0,0,0,
-- M
1,0,0,1,0,
1,1,1,1,0,
1,1,1,1,0,
1,0,0,1,0,
1,0,0,1,0,
1,0,0,1,0,
0,0,0,0,0,
0,0,0,0,0,
-- N
1,0,0,1,0,
1,1,0,1,0,
1,1,0,1,0,
1,0,1,1,0,
1,0,1,1,0,
1,0,0,1,0,
0,0,0,0,0,
0,0,0,0,0,
-- O
0,1,1,0,0,
1,0,0,1,0,
1,0,0,1,0,
1,0,0,1,0,
1,0,0,1,0,
0,1,1,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- P
1,1,1,0,0,
1,0,0,1,0,
1,0,0,1,0,
1,1,1,0,0,
1,0,0,0,0,
1,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- Q
0,1,1,0,0,
1,0,0,1,0,
1,0,0,1,0,
1,0,0,1,0,
1,0,1,1,0,
0,1,1,1,0,
0,0,0,0,0,
0,0,0,0,0,
-- R
1,1,1,0,0,
1,0,0,1,0,
1,1,1,0,0,
1,1,0,0,0,
1,0,1,0,0,
1,0,0,1,0,
0,0,0,0,0,
0,0,0,0,0,
-- S
0,1,1,1,0,
1,0,0,0,0,
0,1,1,0,0,
0,0,0,1,0,
1,0,0,1,0,
0,1,1,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- T
1,1,1,1,1,
0,0,1,0,0,
0,0,1,0,0,
0,0,1,0,0,
0,0,1,0,0,
0,0,1,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- U
1,0,0,1,0,
1,0,0,1,0,
1,0,0,1,0,
1,0,0,1,0,
1,0,0,1,0,
0,1,1,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- V
1,0,0,1,0,
1,0,0,1,0,
1,0,0,1,0,
1,0,0,1,0,
0,1,1,0,0,
0,1,1,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- W
1,0,0,1,0,
1,0,0,1,0,
1,0,0,1,0,
1,0,0,1,0,
1,1,1,1,0,
1,1,1,1,0,
0,0,0,0,0,
0,0,0,0,0,
-- X
1,0,0,1,0,
1,0,0,1,0,
0,1,1,0,0,
0,1,1,0,0,
1,0,0,1,0,
1,0,0,1,0,
0,0,0,0,0,
0,0,0,0,0,
-- Y
1,0,0,0,1,
0,1,0,1,0,
0,1,0,1,0,
0,0,1,0,0,
0,0,1,0,0,
0,0,1,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- Z
1,1,1,1,0,
0,0,0,1,0,
0,0,1,0,0,
0,1,0,0,0,
1,0,0,0,0,
1,1,1,1,0,
0,0,0,0,0,
0,0,0,0,0,
-- [
0,1,1,1,0,
0,1,0,0,0,
0,1,0,0,0,
0,1,0,0,0,
0,1,0,0,0,
0,1,1,1,0,
0,0,0,0,0,
0,0,0,0,0,
-- \
1,0,0,0,0,
0,1,0,0,0,
0,1,0,0,0,
0,0,1,0,0,
0,0,1,0,0,
0,0,0,1,0,
0,0,0,0,0,
0,0,0,0,0,
-- ]
0,1,1,1,0,
0,0,0,1,0,
0,0,0,1,0,
0,0,0,1,0,
0,0,0,1,0,
0,1,1,1,0,
0,0,0,0,0,
0,0,0,0,0,
--       
0,0,1,0,0,
0,1,0,1,0,
0,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
-- _
0,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
0,0,0,0,0,
1,1,1,1,0,
0,0,0,0,0,
0,0,0,0,0,
--
others => 0
);
end package chars;

