package init_message_pkg is

    constant init_message : string := " Z1013.64  v2018.02, 2018-01-30 19:43";
    constant version      : string := "v2018.02";

end package init_message_pkg;
